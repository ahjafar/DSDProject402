// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION
`include "global.v"


module bias_conv1_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV1-1][0:`OUTPUT_NUM_CONV1-1][`WD_BIAS:0] weight	 = {	
		-24'd33091,  -24'd345382,  -24'd986031,  -24'd314271,  24'd400309,  -24'd448129
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_conv1_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV1*`KERNEL_SIZE_CONV1-1][0:`OUTPUT_NUM_CONV1-1][13:0] weight	 = {
14'd247,  14'd464,  -14'd911,  14'd888,  -14'd1589,  -14'd3068,  
14'd950,  -14'd762,  -14'd516,  -14'd343,  -14'd1972,  -14'd1880,  
-14'd1947,  -14'd1365,  -14'd369,  14'd514,  -14'd2763,  14'd71,  
-14'd1916,  -14'd375,  14'd914,  14'd1064,  -14'd2151,  14'd856,  
-14'd3137,  14'd1011,  14'd247,  -14'd666,  -14'd2258,  14'd2362,  

14'd1689,  -14'd776,  -14'd1291,  14'd2099,  -14'd178,  -14'd2206,  
14'd208,  -14'd1154,  -14'd419,  14'd1025,  -14'd2942,  14'd711,  
14'd925,  14'd100,  14'd1016,  14'd1399,  -14'd1774,  14'd1301,  
-14'd1242,  14'd962,  14'd1580,  14'd1905,  -14'd996,  14'd2124,  
-14'd2791,  14'd2,  14'd622,  -14'd1330,  -14'd1809,  -14'd671,  

14'd886,  -14'd385,  -14'd1695,  14'd1718,  14'd355,  -14'd833,  
14'd2550,  14'd212,  14'd987,  14'd888,  14'd744,  14'd711,  
14'd2562,  -14'd257,  14'd1429,  14'd1352,  14'd417,  14'd2049,  
14'd776,  14'd1755,  14'd1958,  14'd1498,  14'd498,  14'd979,  
14'd1253,  14'd1118,  -14'd583,  14'd318,  14'd1914,  -14'd2072,  

-14'd1735,  -14'd378,  -14'd207,  -14'd7,  14'd2647,  14'd163,  
14'd1468,  14'd350,  14'd525,  14'd1304,  14'd2542,  14'd1038,  
14'd75,  14'd2243,  14'd2981,  14'd1678,  14'd1935,  14'd1768,  
14'd2124,  14'd2020,  14'd168,  14'd2411,  14'd2303,  -14'd108,  
14'd720,  -14'd590,  -14'd1400,  14'd2309,  14'd1244,  -14'd3580,  

-14'd1524,  14'd82,  14'd1863,  14'd6,  14'd1707,  14'd442,  
-14'd1060,  14'd1109,  14'd1444,  -14'd1780,  14'd465,  14'd33,  
-14'd735,  14'd53,  14'd1335,  -14'd19,  14'd1379,  14'd1227,  
14'd1149,  14'd2050,  -14'd832,  14'd400,  -14'd222,  -14'd217,  
-14'd442,  14'd1463,  -14'd1258,  14'd1970,  14'd434,  -14'd1883
		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule	


module bias_conv2_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV2-1][0:`OUTPUT_NUM_CONV2-1][`WD_BIAS:0] weight	 = {
	-24'd492928,  -24'd252352,  24'd425549,  -24'd126681,  -24'd362367,  -24'd84127,  24'd122339,  -24'd193094,  24'd178645,  24'd56283,  -24'd15047,  -24'd647019,  -24'd375850,  24'd168062,  -24'd242871,  -24'd1026233		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule



module wieght_conv2_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][`WD:0] weight	 = {
14'd935,  -14'd520,  14'd1060,  14'd504,  -14'd313,  14'd1054,  
-14'd1423,  -14'd1068,  14'd814,  14'd456,  -14'd886,  -14'd1079,  
14'd1276,  -14'd1408,  -14'd1957,  -14'd1050,  -14'd12,  14'd428,  
-14'd59,  14'd403,  -14'd1476,  -14'd499,  -14'd818,  -14'd2231,  
14'd473,  -14'd1360,  -14'd453,  -14'd1395,  -14'd1244,  14'd244,  
-14'd1452,  -14'd830,  14'd562,  -14'd223,  -14'd794,  14'd857,  
14'd272,  14'd349,  -14'd823,  14'd1001,  -14'd636,  14'd252,  
14'd126,  14'd57,  -14'd1241,  14'd270,  -14'd1392,  14'd298,  
14'd245,  -14'd2164,  -14'd1244,  -14'd613,  14'd775,  -14'd984,  
14'd1480,  -14'd1973,  -14'd1964,  -14'd27,  -14'd2855,  14'd1097,  
-14'd1071,  -14'd640,  -14'd76,  -14'd302,  -14'd120,  -14'd2186,  
-14'd717,  -14'd587,  -14'd1290,  -14'd6,  14'd459,  14'd368,  
-14'd435,  -14'd892,  -14'd438,  -14'd492,  14'd225,  14'd827,  
14'd1201,  14'd263,  -14'd629,  14'd1859,  14'd126,  -14'd281,  
14'd120,  14'd919,  -14'd578,  14'd565,  14'd1203,  -14'd1334,  
-14'd685,  14'd485,  -14'd314,  -14'd296,  -14'd714,  -14'd39,  

-14'd560,  14'd45,  -14'd1014,  -14'd1527,  -14'd457,  -14'd638,  
14'd546,  -14'd563,  -14'd619,  14'd1415,  -14'd859,  -14'd931,  
-14'd2687,  -14'd1476,  -14'd49,  -14'd1519,  -14'd769,  -14'd510,  
14'd342,  14'd114,  -14'd591,  -14'd1124,  -14'd125,  14'd535,  
-14'd2066,  -14'd251,  14'd890,  -14'd367,  -14'd1146,  14'd829,  
-14'd325,  14'd1085,  -14'd534,  14'd147,  -14'd292,  -14'd1449,  
-14'd1160,  14'd1096,  -14'd462,  14'd1415,  -14'd205,  14'd1190,  
-14'd569,  -14'd590,  -14'd1032,  14'd687,  -14'd51,  14'd242,  
-14'd544,  -14'd389,  14'd305,  -14'd1090,  14'd65,  -14'd1037,  
-14'd80,  -14'd2025,  14'd1208,  -14'd56,  -14'd1981,  14'd308,  
-14'd451,  -14'd823,  14'd542,  -14'd540,  14'd1755,  14'd117,  
-14'd1763,  -14'd23,  -14'd1477,  14'd688,  14'd510,  -14'd70,  
14'd1022,  -14'd184,  14'd484,  -14'd1568,  -14'd226,  -14'd1429,  
-14'd133,  -14'd1633,  14'd1264,  -14'd104,  14'd1301,  -14'd115,  
14'd662,  14'd388,  14'd1388,  -14'd62,  14'd466,  -14'd1318,  
-14'd583,  14'd977,  -14'd307,  -14'd252,  14'd85,  -14'd925,  

-14'd34,  -14'd467,  14'd185,  -14'd1491,  -14'd268,  -14'd1190,  
14'd1340,  -14'd1197,  -14'd991,  14'd474,  -14'd323,  14'd200,  
-14'd1038,  -14'd463,  -14'd1208,  14'd1599,  -14'd1775,  -14'd1202,  
14'd633,  -14'd230,  14'd567,  -14'd830,  -14'd51,  14'd1422,  
-14'd538,  -14'd834,  14'd234,  14'd174,  -14'd2867,  -14'd526,  
14'd1230,  14'd633,  14'd108,  14'd354,  -14'd317,  -14'd1799,  
14'd296,  -14'd1156,  -14'd58,  -14'd1103,  14'd1195,  14'd489,  
-14'd761,  14'd965,  14'd1210,  14'd309,  -14'd1163,  14'd701,  
-14'd1165,  -14'd208,  -14'd1215,  -14'd787,  -14'd1014,  -14'd1165,  
-14'd286,  -14'd1614,  -14'd950,  -14'd737,  -14'd2465,  14'd813,  
14'd577,  14'd339,  -14'd692,  -14'd641,  14'd958,  -14'd1840,  
14'd1244,  -14'd983,  -14'd1042,  14'd639,  14'd1597,  -14'd876,  
-14'd1259,  -14'd289,  -14'd1100,  -14'd594,  -14'd21,  -14'd207,  
-14'd524,  -14'd470,  -14'd623,  -14'd601,  -14'd1159,  -14'd1233,  
-14'd118,  14'd1153,  -14'd567,  14'd293,  14'd2396,  -14'd785,  
-14'd5,  14'd341,  -14'd60,  14'd1144,  14'd714,  -14'd2911,  

14'd2403,  -14'd992,  -14'd1380,  -14'd304,  -14'd904,  -14'd1978,  
14'd451,  14'd1352,  -14'd795,  14'd919,  -14'd592,  -14'd690,  
14'd663,  14'd295,  14'd961,  14'd394,  -14'd1956,  14'd581,  
-14'd1414,  -14'd1642,  -14'd614,  -14'd1674,  -14'd813,  14'd1286,  
14'd878,  14'd157,  -14'd988,  14'd662,  -14'd2553,  -14'd2060,  
14'd507,  -14'd431,  -14'd299,  -14'd888,  14'd1367,  -14'd1670,  
-14'd746,  -14'd200,  -14'd372,  14'd513,  14'd624,  14'd1030,  
14'd127,  -14'd597,  -14'd468,  14'd54,  -14'd430,  14'd1314,  
-14'd38,  -14'd21,  -14'd139,  -14'd2035,  14'd1012,  14'd692,  
-14'd366,  -14'd388,  14'd1156,  -14'd1199,  -14'd2421,  -14'd391,  
-14'd457,  14'd460,  14'd1197,  -14'd156,  14'd635,  14'd271,  
14'd367,  -14'd859,  -14'd1062,  14'd1399,  -14'd350,  -14'd2515,  
-14'd1077,  14'd295,  14'd627,  -14'd854,  -14'd46,  14'd64,  
-14'd1958,  -14'd69,  -14'd456,  -14'd787,  -14'd2166,  -14'd1154,  
-14'd251,  -14'd1363,  -14'd418,  -14'd887,  14'd765,  -14'd952,  
14'd581,  14'd1524,  -14'd870,  -14'd481,  14'd1823,  -14'd667,  

14'd1349,  -14'd52,  14'd669,  -14'd56,  14'd71,  14'd1065,  
14'd1418,  14'd209,  14'd104,  -14'd680,  14'd1893,  -14'd54,  
-14'd173,  -14'd1047,  14'd433,  14'd367,  -14'd748,  14'd920,  
-14'd783,  -14'd239,  14'd359,  -14'd1001,  14'd84,  14'd1193,  
14'd2156,  14'd673,  -14'd541,  14'd2666,  14'd1702,  14'd329,  
-14'd453,  -14'd956,  -14'd611,  -14'd3018,  -14'd600,  14'd1079,  
-14'd1457,  -14'd1230,  -14'd662,  14'd1074,  -14'd447,  14'd2293,  
14'd277,  -14'd152,  -14'd852,  14'd233,  -14'd1029,  -14'd155,  
-14'd616,  14'd934,  -14'd261,  -14'd852,  14'd558,  -14'd390,  
-14'd1327,  14'd1066,  14'd926,  14'd1362,  -14'd859,  -14'd942,  
-14'd887,  14'd411,  14'd648,  14'd441,  -14'd880,  -14'd288,  
14'd1430,  -14'd1176,  -14'd1962,  -14'd1590,  14'd585,  -14'd2840,  
-14'd187,  14'd732,  14'd958,  14'd773,  -14'd897,  -14'd416,  
14'd1330,  14'd1239,  14'd1735,  -14'd610,  -14'd1825,  14'd1948,  
-14'd397,  -14'd1038,  14'd60,  -14'd715,  14'd1393,  14'd126,  
-14'd305,  14'd379,  14'd330,  14'd77,  14'd1336,  -14'd721,  


-14'd688,  14'd39,  14'd28,  -14'd1360,  14'd41,  -14'd370,  
-14'd91,  -14'd852,  -14'd1423,  -14'd1603,  -14'd1929,  -14'd1441,  
14'd490,  -14'd596,  -14'd3,  -14'd962,  14'd1278,  14'd256,  
-14'd846,  -14'd324,  -14'd1352,  14'd349,  14'd274,  -14'd144,  
14'd1076,  14'd97,  14'd434,  14'd424,  14'd829,  14'd1481,  
-14'd438,  -14'd428,  -14'd984,  -14'd744,  -14'd298,  -14'd362,  
14'd224,  14'd43,  -14'd787,  -14'd338,  -14'd239,  -14'd612,  
14'd1261,  14'd1555,  -14'd655,  14'd864,  -14'd1028,  -14'd1131,  
-14'd659,  14'd91,  -14'd1301,  -14'd1157,  14'd372,  -14'd2609,  
-14'd1087,  -14'd837,  -14'd1568,  -14'd2092,  -14'd863,  14'd27,  
14'd82,  14'd1394,  -14'd896,  14'd987,  14'd535,  -14'd993,  
-14'd479,  -14'd1663,  -14'd429,  -14'd1612,  14'd449,  14'd1594,  
-14'd14,  14'd208,  -14'd305,  -14'd1134,  -14'd1048,  -14'd42,  
-14'd414,  14'd573,  14'd1723,  14'd653,  14'd238,  14'd1050,  
-14'd854,  -14'd907,  -14'd658,  14'd62,  -14'd1152,  -14'd180,  
-14'd243,  -14'd1036,  14'd1149,  14'd525,  14'd994,  14'd631,  

14'd210,  14'd228,  -14'd764,  -14'd821,  -14'd1343,  -14'd1686,  
-14'd325,  14'd712,  14'd608,  14'd504,  -14'd1364,  -14'd578,  
-14'd967,  -14'd857,  -14'd1872,  -14'd376,  14'd120,  -14'd2653,  
14'd468,  14'd534,  14'd782,  14'd749,  -14'd365,  14'd416,  
14'd698,  -14'd700,  14'd1479,  -14'd432,  14'd906,  14'd759,  
14'd712,  -14'd277,  14'd100,  14'd1094,  -14'd1480,  14'd376,  
-14'd129,  14'd371,  14'd1965,  14'd318,  -14'd771,  -14'd191,  
14'd156,  -14'd1062,  14'd400,  14'd749,  -14'd1476,  -14'd660,  
14'd903,  14'd705,  14'd110,  -14'd1029,  14'd206,  14'd706,  
-14'd495,  -14'd370,  -14'd1796,  -14'd689,  -14'd1000,  -14'd2922,  
14'd495,  14'd46,  14'd91,  14'd454,  14'd627,  -14'd1192,  
14'd273,  -14'd89,  14'd384,  -14'd40,  -14'd309,  14'd1046,  
-14'd615,  14'd1211,  14'd1241,  14'd162,  14'd49,  14'd900,  
14'd83,  -14'd543,  14'd962,  -14'd1181,  14'd279,  14'd982,  
-14'd796,  14'd235,  14'd85,  14'd146,  -14'd458,  -14'd660,  
14'd1403,  14'd1355,  14'd407,  14'd104,  14'd1889,  -14'd1290,  

14'd568,  14'd1819,  -14'd654,  14'd483,  -14'd441,  -14'd2127,  
14'd808,  -14'd155,  14'd224,  14'd554,  -14'd1479,  -14'd243,  
-14'd1287,  14'd1017,  -14'd3,  14'd89,  -14'd1895,  -14'd1427,  
14'd1382,  14'd216,  -14'd45,  14'd1033,  -14'd599,  -14'd450,  
-14'd266,  14'd84,  14'd331,  -14'd1671,  14'd1233,  14'd1391,  
14'd1060,  14'd128,  14'd1115,  14'd195,  14'd348,  -14'd1506,  
14'd138,  14'd186,  14'd554,  -14'd97,  14'd29,  14'd924,  
14'd141,  -14'd239,  14'd1606,  14'd535,  -14'd3017,  14'd12,  
-14'd223,  14'd267,  14'd858,  -14'd22,  14'd1544,  14'd996,  
-14'd1419,  14'd286,  -14'd569,  -14'd178,  14'd1704,  14'd1440,  
14'd934,  14'd169,  14'd191,  14'd1161,  14'd1037,  -14'd993,  
14'd509,  14'd857,  -14'd1378,  -14'd1010,  14'd1245,  14'd996,  
-14'd1236,  14'd980,  -14'd127,  14'd832,  14'd628,  14'd424,  
-14'd588,  -14'd938,  -14'd1299,  -14'd1062,  -14'd813,  -14'd797,  
-14'd158,  14'd1328,  -14'd366,  14'd1003,  -14'd1285,  14'd175,  
14'd1459,  14'd494,  14'd1038,  14'd1236,  14'd2726,  -14'd724,  

-14'd65,  -14'd262,  14'd1544,  -14'd223,  -14'd620,  14'd802,  
14'd2037,  14'd813,  14'd340,  14'd661,  -14'd1012,  14'd1764,  
14'd1681,  14'd2031,  14'd140,  14'd148,  -14'd807,  14'd1955,  
14'd205,  14'd1432,  14'd149,  14'd414,  -14'd809,  14'd1293,  
-14'd523,  -14'd1000,  14'd462,  -14'd893,  -14'd54,  14'd717,  
14'd1208,  -14'd324,  -14'd1002,  14'd1051,  14'd127,  -14'd354,  
-14'd355,  14'd220,  14'd1147,  -14'd910,  -14'd1484,  14'd1018,  
14'd131,  -14'd985,  14'd550,  14'd881,  -14'd1643,  14'd930,  
-14'd633,  14'd1302,  -14'd934,  14'd726,  14'd885,  -14'd1632,  
-14'd740,  14'd1221,  14'd1023,  14'd105,  -14'd584,  14'd1339,  
14'd1571,  14'd642,  14'd727,  14'd189,  14'd2430,  -14'd83,  
14'd56,  14'd439,  -14'd280,  14'd716,  -14'd362,  -14'd1095,  
14'd668,  -14'd787,  14'd966,  -14'd1190,  -14'd66,  -14'd410,  
14'd440,  -14'd45,  14'd288,  -14'd954,  -14'd1952,  14'd41,  
-14'd62,  -14'd360,  -14'd175,  14'd66,  -14'd1197,  -14'd197,  
-14'd385,  14'd649,  -14'd559,  14'd1414,  14'd1280,  14'd95,  

14'd490,  -14'd1008,  14'd1941,  14'd1273,  -14'd1138,  14'd1629,  
14'd715,  -14'd1024,  14'd233,  -14'd120,  14'd619,  14'd1001,  
14'd908,  -14'd1693,  14'd154,  14'd552,  -14'd1475,  14'd1184,  
-14'd144,  -14'd727,  14'd329,  14'd378,  -14'd333,  14'd937,  
14'd447,  -14'd853,  -14'd1103,  14'd1064,  -14'd2893,  -14'd1919,  
14'd57,  -14'd219,  14'd973,  14'd141,  -14'd616,  14'd1217,  
-14'd870,  -14'd864,  -14'd978,  -14'd809,  -14'd2888,  14'd304,  
14'd148,  14'd1185,  14'd652,  14'd275,  -14'd152,  -14'd330,  
-14'd513,  -14'd277,  14'd707,  14'd149,  14'd1279,  14'd155,  
-14'd336,  -14'd423,  14'd793,  14'd886,  14'd200,  14'd1294,  
14'd457,  14'd1721,  14'd1795,  -14'd812,  14'd1300,  14'd1452,  
14'd1383,  -14'd1325,  14'd16,  -14'd23,  -14'd1637,  -14'd231,  
-14'd526,  -14'd648,  -14'd74,  14'd807,  14'd139,  14'd781,  
14'd749,  14'd248,  14'd351,  14'd839,  -14'd2612,  14'd894,  
14'd71,  14'd743,  14'd389,  14'd387,  14'd366,  14'd363,  
14'd615,  -14'd2326,  -14'd367,  14'd614,  -14'd68,  -14'd1314,  


-14'd346,  -14'd1273,  -14'd1196,  14'd586,  14'd147,  -14'd2509,  
14'd542,  -14'd355,  14'd195,  14'd629,  -14'd513,  -14'd1828,  
14'd175,  14'd983,  -14'd94,  14'd1777,  14'd1415,  -14'd1958,  
-14'd435,  14'd44,  -14'd1367,  14'd160,  -14'd1283,  -14'd1348,  
14'd534,  -14'd429,  -14'd222,  14'd1359,  14'd902,  14'd1657,  
14'd1822,  14'd590,  -14'd900,  -14'd164,  14'd1481,  -14'd654,  
-14'd1183,  14'd1294,  14'd844,  14'd382,  14'd149,  -14'd948,  
-14'd1405,  -14'd92,  14'd748,  14'd835,  -14'd30,  14'd435,  
14'd802,  14'd1970,  -14'd1733,  -14'd587,  -14'd194,  -14'd161,  
-14'd669,  14'd314,  -14'd48,  -14'd1191,  14'd1529,  -14'd425,  
14'd611,  -14'd585,  14'd14,  14'd1396,  -14'd1691,  -14'd735,  
14'd1058,  -14'd129,  14'd95,  14'd863,  14'd1857,  14'd559,  
14'd6,  14'd1674,  14'd1466,  14'd1073,  14'd627,  14'd529,  
14'd224,  14'd900,  14'd206,  14'd1562,  -14'd189,  14'd1386,  
-14'd1050,  -14'd1652,  14'd293,  14'd610,  -14'd2824,  14'd1126,  
14'd120,  -14'd55,  14'd584,  14'd695,  14'd262,  14'd1208,  

-14'd127,  14'd1121,  14'd296,  14'd198,  14'd1025,  -14'd1627,  
-14'd1293,  14'd300,  14'd1692,  -14'd876,  -14'd91,  14'd2402,  
-14'd2192,  -14'd190,  -14'd260,  -14'd840,  -14'd691,  -14'd251,  
14'd964,  14'd267,  -14'd201,  14'd2223,  -14'd129,  -14'd1082,  
14'd1613,  14'd171,  14'd331,  -14'd869,  14'd495,  14'd705,  
-14'd1796,  -14'd316,  -14'd1009,  14'd1422,  14'd414,  14'd703,  
14'd393,  14'd1426,  14'd1275,  -14'd133,  -14'd2543,  14'd1316,  
14'd229,  -14'd143,  -14'd1538,  14'd1846,  -14'd648,  -14'd815,  
-14'd1015,  -14'd32,  14'd1369,  -14'd1662,  -14'd609,  -14'd67,  
-14'd126,  14'd774,  14'd1185,  -14'd322,  14'd2060,  -14'd829,  
-14'd46,  -14'd52,  -14'd651,  14'd723,  -14'd664,  -14'd50,  
14'd540,  14'd882,  -14'd974,  14'd292,  14'd1242,  14'd389,  
-14'd564,  -14'd698,  14'd824,  14'd1719,  14'd285,  14'd771,  
14'd415,  14'd527,  14'd575,  -14'd1301,  14'd1042,  14'd882,  
-14'd1037,  14'd674,  -14'd1352,  14'd445,  -14'd1394,  -14'd845,  
14'd869,  -14'd508,  14'd367,  -14'd1068,  14'd345,  14'd1214,  

-14'd650,  14'd644,  14'd359,  14'd227,  14'd859,  -14'd134,  
-14'd1249,  -14'd677,  -14'd23,  -14'd714,  -14'd55,  14'd2231,  
-14'd1010,  14'd453,  -14'd553,  14'd436,  -14'd1106,  -14'd791,  
14'd1192,  14'd69,  14'd833,  14'd965,  14'd517,  -14'd2353,  
14'd1241,  -14'd1158,  -14'd611,  14'd501,  14'd271,  14'd400,  
-14'd1570,  14'd249,  14'd542,  14'd1105,  -14'd796,  -14'd1372,  
14'd921,  -14'd885,  14'd2165,  14'd256,  -14'd1482,  14'd932,  
14'd852,  14'd27,  -14'd1067,  14'd1265,  -14'd1386,  -14'd561,  
-14'd263,  -14'd1276,  -14'd802,  -14'd694,  -14'd1265,  14'd551,  
14'd31,  -14'd22,  14'd519,  -14'd29,  14'd1075,  -14'd234,  
14'd624,  14'd861,  -14'd964,  14'd1047,  14'd792,  14'd692,  
14'd877,  14'd475,  -14'd532,  -14'd37,  -14'd995,  14'd781,  
14'd1265,  14'd830,  -14'd483,  14'd1374,  14'd233,  14'd135,  
-14'd1363,  14'd195,  -14'd1135,  -14'd213,  -14'd1997,  -14'd1306,  
14'd1052,  14'd2368,  14'd349,  14'd596,  -14'd2485,  14'd599,  
14'd631,  -14'd1622,  14'd560,  14'd191,  14'd34,  14'd1161,  

-14'd2297,  14'd2123,  14'd2066,  14'd994,  -14'd1334,  14'd2226,  
14'd209,  -14'd900,  -14'd914,  -14'd265,  -14'd2081,  14'd595,  
14'd138,  14'd1130,  14'd1047,  14'd2217,  -14'd2635,  14'd581,  
14'd1207,  14'd835,  14'd278,  14'd1619,  14'd1892,  -14'd1230,  
-14'd1054,  14'd187,  -14'd954,  -14'd1581,  14'd1417,  14'd1625,  
14'd1516,  14'd1519,  14'd612,  14'd897,  -14'd779,  -14'd2057,  
14'd276,  -14'd2214,  -14'd368,  -14'd242,  -14'd979,  14'd746,  
14'd308,  14'd815,  14'd598,  14'd1509,  14'd1452,  14'd261,  
14'd906,  -14'd258,  -14'd925,  -14'd135,  14'd1609,  14'd110,  
14'd1375,  -14'd945,  -14'd1263,  14'd1396,  14'd120,  -14'd2551,  
14'd987,  -14'd1435,  14'd829,  14'd390,  14'd865,  14'd1594,  
14'd517,  14'd167,  14'd1143,  -14'd653,  -14'd980,  14'd820,  
14'd1771,  14'd371,  14'd521,  14'd1638,  14'd230,  -14'd706,  
-14'd1803,  14'd321,  -14'd444,  14'd1097,  -14'd2385,  14'd1889,  
14'd1747,  14'd81,  14'd1514,  -14'd198,  -14'd31,  -14'd1685,  
14'd1139,  -14'd671,  14'd601,  -14'd755,  -14'd1132,  -14'd2113,  

14'd1532,  -14'd534,  14'd785,  14'd291,  -14'd3174,  14'd2602,  
14'd5,  -14'd130,  -14'd1057,  14'd413,  -14'd797,  14'd900,  
14'd881,  14'd146,  -14'd880,  -14'd142,  -14'd2122,  14'd61,  
14'd1250,  14'd1732,  14'd1087,  14'd279,  14'd1593,  14'd380,  
-14'd531,  -14'd389,  -14'd96,  -14'd1079,  14'd543,  14'd1246,  
14'd868,  14'd771,  -14'd428,  14'd1789,  -14'd1198,  14'd120,  
14'd483,  14'd609,  -14'd2369,  -14'd1413,  -14'd2259,  -14'd1888,  
14'd421,  14'd1317,  -14'd1062,  14'd1801,  14'd743,  14'd347,  
14'd1176,  14'd1163,  -14'd997,  14'd755,  14'd1143,  14'd384,  
14'd2054,  -14'd636,  -14'd87,  14'd523,  14'd1086,  -14'd1121,  
14'd84,  -14'd1126,  14'd544,  -14'd1058,  -14'd2937,  14'd1216,  
-14'd969,  14'd951,  14'd2742,  -14'd1539,  -14'd803,  14'd3514,  
14'd204,  14'd726,  14'd1171,  14'd303,  14'd830,  14'd542,  
-14'd189,  14'd1109,  14'd584,  14'd1706,  -14'd2341,  14'd935,  
-14'd107,  14'd344,  14'd29,  14'd22,  14'd183,  -14'd1316,  
14'd1747,  -14'd213,  14'd343,  -14'd637,  -14'd1338,  14'd698,  


14'd1000,  14'd943,  14'd132,  -14'd288,  14'd1729,  -14'd931,  
-14'd189,  14'd711,  14'd953,  -14'd768,  -14'd90,  14'd1181,  
14'd1221,  14'd1468,  14'd844,  14'd708,  14'd1245,  -14'd1676,  
14'd214,  14'd570,  14'd972,  14'd1590,  14'd685,  -14'd1023,  
-14'd1600,  -14'd1262,  14'd353,  -14'd401,  -14'd1928,  14'd187,  
14'd630,  14'd1019,  -14'd684,  14'd1437,  -14'd60,  14'd250,  
-14'd2310,  14'd1170,  14'd1976,  14'd1278,  -14'd1489,  14'd316,  
-14'd228,  -14'd1206,  14'd797,  14'd638,  -14'd1366,  14'd579,  
14'd434,  14'd1614,  14'd1652,  14'd170,  -14'd921,  14'd2619,  
14'd1331,  14'd1125,  -14'd1363,  -14'd177,  14'd1035,  14'd499,  
-14'd1973,  -14'd57,  -14'd1335,  14'd1386,  -14'd1423,  14'd869,  
-14'd145,  -14'd841,  -14'd1028,  14'd24,  14'd807,  14'd689,  
-14'd369,  -14'd749,  14'd95,  14'd1325,  14'd526,  14'd957,  
-14'd243,  14'd132,  -14'd539,  -14'd335,  -14'd224,  14'd199,  
14'd859,  -14'd1284,  14'd399,  -14'd844,  -14'd1792,  -14'd118,  
14'd148,  -14'd832,  -14'd1063,  -14'd666,  -14'd715,  -14'd63,  

-14'd1593,  14'd1625,  14'd1572,  14'd218,  14'd812,  14'd1673,  
-14'd1161,  14'd1071,  14'd2666,  -14'd453,  -14'd1011,  14'd1343,  
14'd417,  -14'd185,  -14'd404,  -14'd111,  14'd598,  -14'd1945,  
14'd400,  -14'd115,  -14'd835,  14'd533,  14'd435,  -14'd927,  
-14'd488,  -14'd163,  14'd107,  14'd50,  14'd82,  14'd116,  
-14'd1933,  14'd506,  14'd652,  14'd414,  -14'd678,  14'd60,  
-14'd71,  -14'd433,  14'd786,  14'd730,  -14'd2005,  -14'd145,  
-14'd1623,  -14'd1047,  -14'd279,  -14'd63,  -14'd3555,  14'd88,  
-14'd1230,  14'd965,  14'd1084,  -14'd920,  -14'd537,  14'd1235,  
14'd37,  14'd879,  14'd718,  14'd1108,  14'd1262,  14'd639,  
-14'd1130,  14'd243,  -14'd253,  -14'd633,  14'd279,  14'd297,  
-14'd299,  14'd527,  14'd236,  -14'd60,  14'd693,  14'd15,  
14'd1938,  -14'd1359,  -14'd560,  -14'd560,  -14'd327,  14'd141,  
14'd438,  14'd575,  14'd767,  -14'd833,  14'd448,  14'd1536,  
14'd1451,  14'd1098,  -14'd1192,  -14'd75,  -14'd1303,  -14'd154,  
14'd395,  -14'd278,  14'd451,  -14'd769,  14'd403,  -14'd610,  

-14'd1724,  -14'd76,  -14'd319,  14'd939,  -14'd1249,  14'd876,  
14'd543,  -14'd1044,  14'd680,  -14'd1725,  -14'd2816,  14'd928,  
-14'd1454,  14'd498,  -14'd635,  14'd246,  -14'd1302,  -14'd1047,  
14'd1017,  14'd469,  -14'd238,  14'd655,  -14'd337,  -14'd1319,  
14'd1128,  14'd305,  14'd1563,  -14'd2,  14'd44,  -14'd100,  
-14'd1828,  -14'd444,  -14'd826,  -14'd1699,  -14'd724,  14'd1733,  
14'd1798,  -14'd837,  -14'd333,  14'd304,  -14'd2343,  14'd194,  
-14'd863,  -14'd1459,  -14'd723,  14'd975,  -14'd1039,  -14'd1492,  
14'd247,  -14'd2439,  -14'd922,  -14'd1047,  -14'd1652,  14'd1009,  
14'd969,  -14'd853,  -14'd400,  -14'd649,  -14'd267,  -14'd1317,  
-14'd999,  -14'd397,  -14'd97,  14'd1103,  14'd1013,  -14'd1533,  
14'd390,  14'd588,  14'd977,  -14'd1056,  14'd827,  14'd537,  
14'd864,  -14'd138,  -14'd1925,  14'd1442,  14'd85,  -14'd426,  
-14'd580,  -14'd936,  -14'd441,  -14'd1366,  -14'd509,  -14'd355,  
14'd278,  14'd1302,  14'd13,  14'd2296,  -14'd1183,  -14'd979,  
-14'd492,  14'd43,  -14'd1112,  -14'd1512,  14'd726,  -14'd1820,  

14'd120,  -14'd433,  -14'd1377,  14'd224,  -14'd4355,  -14'd1039,  
-14'd686,  -14'd726,  -14'd1530,  -14'd342,  -14'd3089,  -14'd692,  
-14'd1068,  14'd8,  14'd809,  14'd822,  -14'd3312,  14'd1073,  
-14'd141,  -14'd744,  -14'd1070,  14'd1434,  14'd1176,  -14'd547,  
14'd719,  14'd1489,  -14'd488,  14'd142,  14'd1718,  -14'd1979,  
14'd924,  -14'd1129,  -14'd757,  14'd735,  -14'd2641,  -14'd642,  
14'd274,  -14'd852,  -14'd2153,  -14'd1493,  -14'd685,  -14'd1782,  
14'd1543,  -14'd245,  -14'd1051,  14'd312,  -14'd613,  -14'd2415,  
14'd2259,  14'd1240,  -14'd924,  -14'd1141,  -14'd406,  -14'd1003,  
-14'd151,  14'd204,  -14'd361,  -14'd153,  14'd486,  -14'd1957,  
-14'd748,  -14'd2625,  -14'd1861,  -14'd958,  -14'd96,  -14'd904,  
-14'd1044,  -14'd392,  14'd917,  14'd1282,  -14'd853,  14'd1031,  
-14'd442,  -14'd878,  -14'd953,  14'd1744,  14'd977,  -14'd2234,  
-14'd977,  14'd81,  14'd382,  14'd67,  -14'd2279,  14'd1286,  
14'd865,  14'd451,  -14'd463,  14'd1487,  14'd650,  -14'd379,  
-14'd1322,  14'd454,  -14'd149,  -14'd359,  -14'd638,  14'd405,  

-14'd362,  14'd182,  -14'd229,  14'd557,  -14'd1476,  14'd513,  
14'd516,  14'd1485,  14'd378,  14'd159,  -14'd1503,  14'd1953,  
14'd1061,  -14'd194,  14'd519,  14'd499,  -14'd914,  -14'd1200,  
14'd2181,  14'd503,  14'd97,  14'd397,  14'd1024,  -14'd520,  
14'd540,  14'd320,  14'd291,  -14'd253,  14'd477,  -14'd566,  
14'd1195,  -14'd101,  14'd482,  14'd1994,  -14'd120,  -14'd1946,  
-14'd88,  14'd1087,  -14'd499,  -14'd1357,  -14'd174,  -14'd98,  
14'd1542,  14'd394,  -14'd295,  14'd1021,  14'd1541,  -14'd2147,  
14'd2485,  -14'd805,  -14'd1864,  -14'd308,  14'd2212,  -14'd65,  
14'd336,  -14'd54,  -14'd1101,  14'd655,  -14'd1581,  -14'd1458,  
-14'd1116,  -14'd918,  -14'd2603,  -14'd2201,  14'd511,  -14'd1247,  
-14'd1217,  14'd136,  -14'd164,  14'd574,  -14'd3331,  14'd2512,  
14'd226,  -14'd190,  -14'd130,  -14'd1002,  14'd1334,  -14'd675,  
14'd1317,  -14'd627,  14'd1536,  14'd1306,  -14'd1870,  14'd276,  
14'd1498,  14'd69,  14'd155,  14'd1368,  -14'd66,  -14'd123,  
14'd24,  -14'd711,  14'd374,  14'd723,  -14'd1436,  14'd1817,  


-14'd503,  14'd51,  -14'd670,  -14'd1902,  14'd1113,  14'd1892,  
-14'd1825,  14'd720,  -14'd208,  -14'd177,  -14'd547,  -14'd131,  
14'd2152,  -14'd713,  -14'd756,  14'd406,  -14'd267,  -14'd611,  
-14'd1421,  -14'd1270,  14'd416,  -14'd158,  -14'd754,  -14'd553,  
14'd674,  14'd564,  -14'd422,  -14'd1441,  14'd162,  -14'd646,  
-14'd1499,  14'd1562,  14'd882,  -14'd347,  -14'd1109,  14'd922,  
-14'd228,  14'd1355,  14'd2209,  14'd324,  -14'd1219,  14'd69,  
-14'd941,  -14'd1551,  14'd911,  14'd271,  14'd881,  -14'd1975,  
-14'd1412,  14'd2656,  14'd3031,  14'd1715,  -14'd3077,  14'd1789,  
14'd1543,  -14'd911,  14'd558,  14'd405,  -14'd609,  14'd99,  
-14'd1160,  14'd775,  14'd328,  -14'd263,  -14'd627,  14'd1132,  
-14'd1323,  14'd575,  -14'd1436,  -14'd309,  -14'd1366,  14'd427,  
14'd453,  -14'd1006,  -14'd2203,  -14'd1649,  14'd705,  -14'd559,  
-14'd274,  14'd1277,  14'd1144,  14'd529,  -14'd1170,  -14'd147,  
-14'd247,  -14'd457,  -14'd680,  -14'd220,  -14'd1641,  -14'd307,  
14'd312,  -14'd499,  -14'd1303,  -14'd1225,  14'd1411,  -14'd20,  

-14'd1121,  14'd393,  14'd1131,  -14'd501,  -14'd1664,  14'd677,  
-14'd1412,  14'd1009,  14'd773,  -14'd349,  -14'd2868,  14'd1568,  
14'd438,  14'd719,  14'd809,  -14'd113,  14'd368,  -14'd1623,  
-14'd630,  -14'd2136,  -14'd460,  14'd357,  -14'd1968,  14'd970,  
-14'd308,  -14'd236,  -14'd130,  -14'd1062,  14'd49,  14'd1907,  
-14'd349,  14'd230,  14'd68,  -14'd258,  -14'd665,  14'd1087,  
14'd1116,  14'd637,  -14'd93,  14'd366,  -14'd2308,  14'd1639,  
-14'd1929,  -14'd295,  -14'd1630,  -14'd845,  -14'd909,  -14'd33,  
14'd1203,  14'd1250,  14'd1851,  14'd1155,  -14'd2931,  14'd2175,  
14'd1719,  14'd237,  -14'd1086,  14'd1065,  14'd973,  -14'd2334,  
14'd386,  -14'd2000,  -14'd1571,  -14'd1087,  14'd2039,  -14'd172,  
-14'd68,  14'd808,  14'd174,  -14'd487,  -14'd575,  -14'd52,  
-14'd55,  -14'd1531,  -14'd772,  -14'd618,  14'd2224,  -14'd694,  
-14'd701,  -14'd276,  14'd1716,  14'd196,  -14'd628,  -14'd119,  
-14'd1261,  14'd271,  -14'd462,  -14'd2075,  -14'd927,  -14'd807,  
14'd971,  14'd339,  -14'd437,  -14'd142,  14'd1562,  -14'd831,  

-14'd1095,  14'd947,  -14'd495,  14'd1052,  -14'd3157,  14'd186,  
14'd1730,  -14'd1677,  -14'd786,  14'd304,  -14'd796,  14'd304,  
-14'd502,  14'd1320,  -14'd933,  14'd88,  -14'd979,  14'd495,  
-14'd924,  -14'd1912,  -14'd1064,  14'd768,  -14'd810,  -14'd991,  
-14'd1244,  14'd773,  14'd626,  -14'd85,  -14'd425,  14'd268,  
-14'd841,  -14'd2427,  14'd335,  -14'd471,  -14'd1180,  14'd301,  
14'd629,  -14'd1488,  -14'd572,  -14'd121,  -14'd1121,  -14'd1068,  
-14'd877,  -14'd916,  14'd703,  -14'd474,  -14'd31,  -14'd452,  
14'd1366,  14'd699,  -14'd762,  14'd442,  -14'd322,  -14'd536,  
14'd897,  14'd1359,  -14'd1214,  -14'd548,  14'd402,  -14'd2162,  
-14'd1422,  14'd288,  -14'd2261,  -14'd1194,  14'd442,  -14'd3179,  
-14'd1570,  14'd28,  14'd614,  14'd1016,  -14'd946,  14'd1941,  
-14'd780,  14'd176,  -14'd975,  -14'd700,  14'd1201,  -14'd132,  
-14'd489,  14'd251,  14'd803,  -14'd685,  14'd1218,  -14'd751,  
-14'd425,  -14'd1134,  -14'd561,  14'd133,  -14'd1549,  -14'd1737,  
-14'd263,  14'd542,  -14'd460,  -14'd1297,  14'd1001,  14'd1953,  

14'd1437,  -14'd960,  -14'd1217,  14'd660,  -14'd1751,  -14'd852,  
-14'd179,  14'd91,  14'd832,  -14'd631,  -14'd623,  14'd741,  
14'd310,  14'd395,  14'd581,  14'd401,  -14'd1851,  14'd1988,  
-14'd1564,  -14'd1997,  -14'd1745,  -14'd405,  -14'd1770,  -14'd1694,  
14'd527,  14'd30,  14'd1191,  -14'd239,  -14'd309,  -14'd458,  
14'd190,  -14'd132,  -14'd709,  -14'd173,  -14'd263,  -14'd1685,  
14'd45,  14'd603,  -14'd986,  14'd370,  14'd1556,  -14'd1504,  
-14'd1269,  -14'd1165,  14'd191,  -14'd1023,  -14'd456,  14'd347,  
-14'd1489,  -14'd171,  -14'd1219,  -14'd1928,  14'd174,  14'd471,  
14'd735,  14'd1175,  -14'd622,  14'd121,  14'd2549,  14'd404,  
-14'd1050,  -14'd1253,  -14'd1613,  -14'd2469,  14'd732,  -14'd1765,  
14'd344,  -14'd2005,  -14'd501,  14'd422,  14'd136,  14'd466,  
-14'd2449,  -14'd720,  -14'd32,  -14'd1858,  -14'd189,  -14'd817,  
14'd476,  14'd1237,  14'd1475,  -14'd25,  -14'd1236,  14'd162,  
14'd1089,  14'd77,  -14'd963,  14'd477,  -14'd827,  -14'd212,  
-14'd1732,  14'd367,  14'd1005,  -14'd384,  -14'd619,  14'd18,  

-14'd288,  -14'd979,  -14'd1956,  14'd924,  -14'd894,  -14'd1442,  
-14'd823,  -14'd57,  14'd1823,  14'd827,  -14'd1161,  14'd1892,  
14'd1384,  -14'd1451,  -14'd1067,  14'd1489,  -14'd544,  14'd127,  
-14'd400,  -14'd931,  -14'd392,  -14'd824,  -14'd931,  -14'd1757,  
14'd451,  -14'd255,  -14'd354,  14'd155,  -14'd167,  -14'd117,  
-14'd166,  -14'd1627,  -14'd974,  -14'd564,  -14'd1827,  -14'd376,  
14'd748,  14'd1976,  -14'd300,  -14'd200,  14'd633,  14'd574,  
-14'd1407,  -14'd866,  -14'd1012,  -14'd553,  -14'd125,  14'd692,  
14'd977,  -14'd1910,  -14'd588,  -14'd531,  14'd37,  -14'd197,  
-14'd10,  -14'd992,  14'd602,  -14'd998,  14'd407,  -14'd1610,  
-14'd1613,  14'd1715,  -14'd432,  -14'd1345,  14'd549,  -14'd1110,  
-14'd191,  -14'd92,  -14'd162,  14'd274,  14'd421,  -14'd2795,  
-14'd2646,  -14'd1201,  14'd263,  -14'd1873,  -14'd1976,  14'd1085,  
14'd1743,  14'd1291,  -14'd340,  14'd208,  -14'd1397,  -14'd317,  
14'd873,  -14'd2006,  14'd434,  -14'd67,  -14'd678,  -14'd578,  
-14'd366,  -14'd436,  -14'd84,  14'd853,  -14'd1274,  14'd199
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule


module bias_fc1_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC1-1][0:`OUTPUT_NUM_FC1-1][`WD_BIAS:0] weight	 = {
-24'd219560,  -24'd253697,  -24'd55433,  -24'd97677,  24'd293697,  -24'd243881,  24'd320084,  24'd224550,  24'd239030,  24'd511222,  24'd91710,  24'd236129,  24'd189478,  24'd189715,  24'd237750,  24'd85050,  
24'd84279,  -24'd41102,  24'd389770,  24'd141391,  -24'd114359,  24'd179309,  24'd335280,  24'd91496,  -24'd304524,  24'd51767,  24'd50531,  24'd398249,  24'd125193,  24'd59246,  24'd302096,  -24'd391546,  
-24'd8719,  -24'd143200,  24'd86710,  -24'd121286,  -24'd17574,  24'd193986,  24'd334251,  24'd418338,  -24'd29725,  -24'd164781,  24'd19566,  24'd369659,  24'd369117,  24'd485986,  24'd255667,  24'd184972,  
-24'd350874,  24'd83616,  -24'd113753,  24'd50318,  -24'd218172,  24'd245365,  -24'd212866,  -24'd167942,  24'd24266,  -24'd290894,  -24'd45370,  24'd333035,  24'd76391,  24'd331919,  24'd249570,  24'd116175,  
24'd314113,  24'd322302,  -24'd387295,  -24'd139803,  24'd555959,  24'd41557,  -24'd71756,  24'd250106,  24'd125286,  24'd209370,  -24'd167080,  24'd330490,  24'd186924,  24'd87729,  -24'd220844,  24'd340936,  
-24'd135930,  24'd117423,  24'd224274,  -24'd3834,  -24'd49645,  -24'd105418,  24'd52762,  24'd96732,  -24'd152523,  24'd141711,  24'd257837,  -24'd91013,  24'd178395,  24'd55568,  -24'd93767,  -24'd131308,  
24'd155983,  -24'd449369,  24'd184192,  -24'd39257,  -24'd140313,  24'd360847,  24'd255272,  24'd73788,  -24'd213748,  24'd163158,  24'd149546,  24'd206663,  -24'd58642,  -24'd77157,  -24'd41775,  24'd140758,  
24'd396969,  24'd190957,  24'd87027,  -24'd48891,  24'd157309,  -24'd282668,  -24'd283377,  -24'd195665
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_fc1_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1*`OUTPUT_BATCH_FC1)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV2*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC1*`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1-1][0:`OUTPUT_NUM_FC1-1][0:`OUTPUT_NUM_CONV2-1][`WD:0] weight	 = {
-14'd353,  14'd196,  -14'd208,  14'd2001,  -14'd16,  14'd3,  14'd483,  -14'd1753,  14'd896,  14'd557,  -14'd283,  -14'd533,  14'd823,  -14'd921,  -14'd713,  -14'd193,  
14'd1758,  14'd186,  14'd961,  14'd846,  -14'd870,  14'd662,  -14'd1155,  14'd980,  14'd170,  -14'd119,  14'd16,  14'd263,  14'd1008,  -14'd562,  -14'd55,  14'd305,  
14'd644,  -14'd1114,  14'd340,  -14'd1010,  -14'd1352,  -14'd622,  14'd171,  -14'd1148,  14'd484,  -14'd940,  14'd1716,  14'd1024,  14'd1260,  -14'd586,  -14'd880,  14'd1980,  
14'd481,  14'd213,  14'd732,  14'd2,  -14'd803,  14'd1339,  14'd1717,  14'd573,  14'd1285,  -14'd32,  14'd1141,  14'd15,  14'd703,  14'd1411,  -14'd444,  -14'd174,  
14'd1834,  14'd1638,  -14'd1313,  14'd641,  14'd1877,  14'd1347,  14'd1297,  14'd1158,  14'd783,  -14'd520,  14'd185,  14'd1319,  14'd1829,  14'd701,  -14'd2033,  14'd528,  
14'd1030,  14'd680,  -14'd1018,  14'd744,  14'd844,  -14'd341,  14'd772,  -14'd1615,  -14'd558,  -14'd803,  14'd2106,  -14'd465,  -14'd137,  -14'd919,  14'd1528,  -14'd53,  
14'd163,  14'd535,  -14'd594,  -14'd675,  -14'd145,  14'd787,  14'd391,  -14'd56,  14'd584,  14'd365,  14'd1731,  14'd486,  -14'd1152,  -14'd604,  -14'd1902,  -14'd1421,  
14'd335,  -14'd1065,  -14'd560,  -14'd895,  -14'd101,  14'd426,  14'd204,  -14'd992,  14'd273,  14'd1396,  -14'd201,  14'd476,  14'd1670,  -14'd194,  -14'd736,  14'd597,  
14'd1126,  -14'd1343,  -14'd960,  -14'd1332,  -14'd87,  14'd253,  -14'd631,  -14'd1234,  -14'd1149,  -14'd1767,  -14'd752,  -14'd682,  14'd1060,  14'd1433,  14'd594,  14'd446,  
-14'd359,  -14'd144,  -14'd3010,  -14'd594,  -14'd834,  -14'd446,  -14'd93,  -14'd200,  -14'd1068,  -14'd1205,  14'd699,  -14'd854,  -14'd731,  -14'd746,  14'd744,  -14'd1290,  
-14'd371,  14'd140,  14'd1647,  -14'd1760,  -14'd447,  -14'd1015,  -14'd197,  -14'd959,  -14'd487,  -14'd1042,  -14'd1229,  14'd553,  14'd647,  -14'd225,  -14'd52,  -14'd161,  
-14'd100,  14'd1351,  14'd886,  -14'd1412,  -14'd1133,  14'd24,  14'd869,  -14'd386,  14'd589,  14'd506,  -14'd1313,  -14'd248,  -14'd1218,  14'd1440,  -14'd1045,  -14'd437,  
-14'd9,  -14'd659,  -14'd896,  -14'd1216,  -14'd822,  -14'd1069,  -14'd1140,  -14'd1434,  -14'd1212,  -14'd703,  -14'd1900,  -14'd820,  14'd353,  14'd1530,  -14'd687,  -14'd532,  
14'd17,  -14'd654,  14'd1228,  14'd785,  -14'd14,  -14'd2633,  -14'd463,  -14'd456,  14'd78,  14'd922,  -14'd1480,  -14'd939,  14'd72,  14'd946,  -14'd1084,  -14'd25,  
-14'd2172,  -14'd1372,  14'd563,  14'd703,  -14'd241,  -14'd1868,  14'd154,  -14'd1521,  -14'd14,  14'd1580,  -14'd114,  14'd806,  -14'd1018,  -14'd450,  -14'd22,  -14'd1996,  
-14'd502,  -14'd665,  14'd270,  14'd1345,  14'd954,  -14'd139,  -14'd2309,  -14'd298,  14'd672,  -14'd28,  -14'd1282,  -14'd1259,  14'd410,  -14'd63,  14'd1809,  -14'd246,  
-14'd865,  -14'd1465,  -14'd288,  14'd2405,  14'd789,  -14'd206,  -14'd648,  14'd744,  -14'd775,  -14'd59,  14'd1665,  -14'd1105,  -14'd157,  -14'd469,  -14'd267,  -14'd1380,  
14'd75,  -14'd209,  14'd447,  14'd185,  -14'd374,  -14'd1602,  -14'd2730,  14'd153,  -14'd2423,  14'd1369,  -14'd220,  -14'd791,  14'd787,  14'd10,  -14'd343,  14'd1362,  
-14'd246,  -14'd972,  14'd466,  14'd734,  -14'd1419,  14'd154,  14'd196,  -14'd60,  -14'd672,  -14'd1337,  -14'd1245,  14'd1374,  14'd1313,  -14'd21,  14'd271,  14'd901,  
-14'd683,  -14'd942,  -14'd754,  -14'd566,  -14'd386,  -14'd225,  14'd1164,  14'd304,  14'd1115,  -14'd970,  14'd143,  14'd1623,  -14'd323,  -14'd299,  -14'd35,  -14'd550,  
-14'd1045,  14'd1470,  -14'd1105,  -14'd825,  14'd216,  14'd577,  -14'd1071,  14'd724,  14'd2756,  14'd374,  14'd2176,  -14'd1596,  -14'd50,  -14'd1335,  14'd132,  -14'd31,  
-14'd843,  14'd308,  -14'd2074,  -14'd768,  -14'd594,  -14'd835,  -14'd2325,  -14'd1334,  14'd1255,  -14'd1487,  14'd786,  14'd89,  -14'd224,  -14'd2315,  14'd106,  14'd1161,  
14'd138,  -14'd203,  -14'd1464,  14'd182,  -14'd2323,  -14'd1112,  -14'd1744,  14'd702,  -14'd677,  -14'd482,  14'd861,  -14'd245,  -14'd469,  14'd1600,  14'd306,  -14'd121,  
-14'd873,  14'd143,  14'd1966,  -14'd1300,  -14'd1472,  -14'd32,  14'd1491,  -14'd881,  14'd37,  -14'd363,  -14'd760,  14'd339,  14'd320,  14'd2347,  14'd1646,  14'd822,  
14'd1330,  14'd456,  14'd1315,  14'd952,  -14'd11,  14'd655,  14'd1344,  14'd261,  14'd240,  -14'd2247,  -14'd698,  14'd841,  -14'd498,  -14'd473,  14'd921,  14'd984,  

-14'd425,  -14'd6,  -14'd265,  14'd480,  -14'd554,  14'd804,  -14'd1110,  -14'd207,  -14'd1525,  -14'd351,  14'd103,  14'd579,  -14'd174,  -14'd414,  14'd412,  14'd749,  
-14'd1250,  -14'd1365,  -14'd755,  -14'd824,  -14'd1224,  -14'd930,  -14'd108,  -14'd216,  14'd112,  -14'd1008,  14'd331,  14'd1067,  14'd1109,  14'd406,  -14'd1746,  -14'd845,  
-14'd456,  -14'd837,  -14'd492,  -14'd692,  -14'd226,  14'd1082,  -14'd472,  14'd687,  14'd435,  -14'd1274,  -14'd421,  -14'd770,  -14'd222,  14'd364,  14'd488,  -14'd920,  
14'd548,  14'd750,  -14'd147,  14'd390,  -14'd512,  -14'd117,  -14'd1703,  -14'd634,  -14'd924,  -14'd312,  -14'd1781,  -14'd226,  -14'd657,  -14'd509,  14'd20,  14'd30,  
14'd1405,  -14'd554,  -14'd341,  -14'd909,  14'd529,  -14'd1704,  -14'd610,  -14'd344,  -14'd715,  14'd445,  -14'd1658,  -14'd79,  14'd336,  14'd278,  -14'd133,  -14'd1559,  
14'd254,  14'd47,  14'd1097,  -14'd822,  14'd352,  14'd744,  -14'd629,  -14'd959,  -14'd454,  14'd959,  -14'd1098,  14'd404,  14'd1413,  14'd139,  -14'd530,  -14'd1548,  
-14'd222,  -14'd401,  -14'd1001,  -14'd315,  -14'd253,  -14'd356,  14'd474,  -14'd704,  -14'd1055,  14'd1068,  14'd640,  -14'd1314,  -14'd43,  14'd489,  -14'd271,  -14'd1074,  
14'd945,  -14'd851,  14'd338,  14'd750,  14'd823,  14'd762,  -14'd1088,  14'd317,  14'd429,  14'd289,  -14'd282,  14'd622,  -14'd379,  -14'd286,  14'd746,  14'd683,  
-14'd42,  -14'd1211,  14'd37,  -14'd939,  -14'd353,  14'd321,  14'd764,  -14'd921,  14'd199,  -14'd162,  -14'd140,  -14'd1064,  -14'd1986,  -14'd780,  14'd44,  -14'd1836,  
14'd209,  -14'd269,  -14'd288,  -14'd794,  14'd371,  14'd127,  -14'd900,  -14'd278,  14'd314,  14'd242,  -14'd38,  -14'd198,  14'd92,  -14'd341,  -14'd1557,  -14'd1181,  
-14'd519,  -14'd508,  -14'd65,  -14'd1577,  -14'd1458,  -14'd365,  -14'd1066,  -14'd18,  -14'd1605,  14'd256,  14'd287,  -14'd607,  -14'd837,  14'd36,  -14'd312,  -14'd75,  
-14'd1629,  -14'd1517,  -14'd72,  -14'd560,  14'd625,  -14'd1101,  14'd142,  -14'd251,  14'd428,  14'd1154,  14'd206,  -14'd797,  14'd434,  -14'd293,  -14'd69,  14'd155,  
14'd208,  14'd88,  -14'd1449,  14'd749,  14'd680,  -14'd1091,  14'd126,  -14'd796,  14'd568,  -14'd679,  14'd515,  14'd1103,  14'd457,  -14'd886,  14'd505,  -14'd932,  
-14'd173,  -14'd290,  -14'd746,  14'd1096,  -14'd1279,  14'd918,  14'd397,  -14'd457,  -14'd508,  -14'd1639,  -14'd943,  -14'd824,  14'd337,  14'd518,  -14'd774,  14'd275,  
-14'd392,  -14'd269,  14'd187,  -14'd816,  14'd761,  -14'd298,  -14'd1362,  14'd596,  -14'd377,  -14'd234,  -14'd558,  -14'd587,  -14'd498,  -14'd636,  -14'd940,  -14'd519,  
14'd1182,  14'd376,  -14'd844,  -14'd840,  -14'd784,  -14'd481,  -14'd1514,  -14'd943,  14'd805,  -14'd855,  -14'd1342,  14'd89,  -14'd100,  -14'd608,  -14'd685,  -14'd766,  
-14'd1617,  14'd539,  -14'd118,  14'd521,  -14'd754,  14'd380,  14'd350,  -14'd227,  -14'd1479,  14'd345,  -14'd589,  -14'd1202,  -14'd1577,  -14'd651,  -14'd1064,  14'd1045,  
14'd269,  14'd964,  14'd43,  14'd754,  14'd1030,  -14'd600,  14'd645,  -14'd620,  -14'd1039,  14'd82,  -14'd753,  14'd990,  -14'd20,  -14'd483,  14'd455,  -14'd1076,  
-14'd156,  -14'd449,  -14'd255,  -14'd643,  -14'd770,  14'd176,  -14'd1019,  -14'd407,  14'd139,  14'd453,  -14'd741,  -14'd1071,  -14'd1401,  -14'd378,  -14'd548,  -14'd724,  
14'd221,  -14'd919,  -14'd58,  -14'd536,  -14'd989,  -14'd871,  -14'd4,  -14'd1533,  -14'd100,  -14'd452,  -14'd1124,  14'd726,  14'd286,  -14'd1173,  14'd393,  14'd40,  
-14'd838,  14'd293,  14'd577,  -14'd982,  -14'd1395,  -14'd184,  -14'd1278,  14'd187,  -14'd60,  -14'd1675,  14'd254,  -14'd370,  -14'd531,  -14'd1697,  14'd471,  14'd97,  
14'd749,  -14'd1419,  -14'd404,  -14'd309,  -14'd655,  -14'd769,  -14'd317,  14'd87,  14'd1194,  -14'd318,  -14'd1588,  14'd15,  14'd783,  -14'd1162,  -14'd67,  -14'd955,  
14'd182,  -14'd137,  14'd1327,  14'd193,  -14'd884,  -14'd389,  14'd913,  14'd249,  14'd278,  14'd965,  14'd187,  -14'd1337,  -14'd628,  -14'd105,  -14'd600,  14'd792,  
-14'd719,  -14'd1293,  14'd192,  -14'd1179,  -14'd205,  14'd916,  -14'd332,  -14'd177,  -14'd496,  -14'd549,  -14'd157,  -14'd164,  -14'd682,  -14'd1043,  14'd462,  -14'd170,  
-14'd317,  -14'd985,  14'd185,  14'd1287,  -14'd530,  -14'd1033,  -14'd1389,  -14'd830,  14'd608,  14'd75,  14'd259,  -14'd255,  -14'd86,  -14'd927,  14'd715,  14'd527,  

-14'd870,  -14'd938,  14'd1563,  -14'd867,  -14'd1003,  14'd522,  -14'd2474,  14'd399,  14'd1241,  -14'd1098,  -14'd1872,  14'd242,  -14'd245,  14'd395,  14'd1218,  14'd207,  
14'd251,  -14'd403,  14'd3065,  -14'd372,  -14'd132,  14'd655,  14'd205,  -14'd1437,  14'd264,  14'd1255,  -14'd2410,  14'd650,  14'd504,  -14'd416,  14'd479,  -14'd728,  
-14'd1053,  14'd131,  14'd284,  -14'd1202,  14'd1067,  14'd341,  14'd1421,  -14'd448,  -14'd516,  14'd61,  -14'd62,  14'd1015,  -14'd813,  14'd3860,  -14'd279,  -14'd809,  
-14'd946,  14'd965,  14'd945,  14'd888,  -14'd176,  14'd121,  14'd959,  -14'd548,  14'd1328,  -14'd44,  -14'd193,  -14'd1163,  -14'd1253,  14'd1904,  14'd535,  -14'd17,  
14'd2013,  14'd2477,  -14'd512,  -14'd449,  -14'd261,  -14'd267,  14'd1660,  14'd655,  14'd702,  14'd191,  -14'd699,  14'd219,  -14'd722,  -14'd741,  14'd370,  14'd825,  
14'd7,  14'd192,  14'd1672,  14'd1301,  14'd1039,  14'd426,  -14'd2316,  14'd637,  -14'd1344,  14'd929,  -14'd1280,  -14'd196,  -14'd465,  14'd1055,  -14'd19,  14'd485,  
-14'd370,  14'd988,  14'd57,  -14'd764,  -14'd200,  -14'd197,  14'd666,  14'd702,  14'd53,  14'd424,  14'd166,  -14'd71,  -14'd64,  -14'd817,  14'd538,  -14'd758,  
-14'd877,  -14'd1898,  14'd951,  -14'd1269,  -14'd1609,  -14'd1197,  14'd657,  14'd318,  14'd27,  -14'd313,  -14'd1626,  -14'd920,  -14'd519,  14'd177,  14'd1435,  -14'd136,  
14'd861,  14'd30,  -14'd198,  -14'd370,  -14'd1203,  14'd4,  14'd68,  -14'd694,  14'd561,  -14'd1086,  -14'd17,  -14'd613,  -14'd105,  14'd1388,  -14'd768,  -14'd1331,  
14'd2194,  14'd542,  -14'd347,  -14'd547,  -14'd416,  -14'd740,  14'd1845,  -14'd482,  14'd1274,  -14'd501,  14'd740,  14'd407,  14'd2155,  14'd813,  -14'd527,  14'd728,  
14'd440,  14'd200,  14'd292,  -14'd619,  14'd1163,  -14'd514,  -14'd640,  14'd215,  -14'd980,  -14'd1200,  14'd0,  14'd491,  -14'd1599,  -14'd22,  -14'd146,  14'd313,  
14'd1003,  14'd1076,  14'd454,  -14'd85,  14'd273,  -14'd94,  -14'd199,  14'd1346,  -14'd1545,  -14'd501,  14'd102,  -14'd707,  -14'd502,  -14'd40,  14'd115,  -14'd510,  
14'd687,  14'd1587,  -14'd1179,  -14'd646,  14'd61,  14'd1503,  14'd202,  14'd459,  14'd911,  14'd792,  14'd377,  -14'd1181,  14'd1496,  -14'd1506,  -14'd1025,  -14'd1664,  
14'd203,  -14'd391,  14'd506,  14'd1813,  14'd380,  14'd912,  -14'd784,  14'd1287,  -14'd409,  -14'd306,  14'd174,  -14'd800,  -14'd85,  14'd413,  14'd374,  -14'd81,  
14'd2631,  14'd1582,  -14'd542,  -14'd228,  14'd469,  14'd513,  -14'd875,  -14'd907,  14'd507,  -14'd1276,  -14'd580,  14'd186,  14'd1928,  -14'd653,  14'd930,  14'd1728,  
14'd1566,  -14'd1128,  -14'd472,  -14'd197,  -14'd1051,  -14'd924,  14'd421,  -14'd983,  14'd42,  -14'd984,  -14'd1445,  14'd1412,  -14'd1644,  14'd204,  -14'd708,  14'd60,  
14'd1633,  14'd968,  14'd852,  -14'd757,  -14'd565,  14'd219,  14'd666,  -14'd324,  14'd1315,  14'd1455,  -14'd1239,  14'd244,  14'd1023,  14'd2259,  -14'd510,  14'd180,  
-14'd543,  -14'd66,  -14'd869,  14'd1262,  14'd537,  -14'd282,  14'd432,  14'd90,  14'd1051,  -14'd87,  14'd841,  14'd222,  -14'd17,  -14'd407,  -14'd1126,  14'd288,  
-14'd1595,  14'd256,  -14'd1612,  -14'd1203,  -14'd24,  -14'd1070,  -14'd191,  14'd1470,  -14'd1749,  14'd1495,  -14'd513,  -14'd512,  -14'd2164,  -14'd550,  -14'd691,  14'd724,  
14'd271,  -14'd1143,  -14'd974,  -14'd1582,  14'd290,  -14'd893,  -14'd561,  -14'd572,  -14'd1155,  -14'd696,  -14'd79,  14'd472,  14'd752,  -14'd245,  -14'd1519,  14'd118,  
14'd2328,  14'd307,  14'd1894,  -14'd821,  -14'd1169,  14'd1343,  -14'd414,  14'd1242,  14'd408,  14'd1473,  -14'd9,  14'd1294,  14'd162,  14'd2311,  14'd1023,  14'd1173,  
14'd214,  -14'd478,  14'd1422,  14'd608,  14'd169,  -14'd1579,  -14'd398,  14'd779,  14'd858,  -14'd664,  14'd324,  14'd1220,  14'd402,  14'd708,  -14'd477,  -14'd686,  
-14'd1095,  14'd265,  -14'd523,  -14'd366,  -14'd273,  -14'd573,  14'd46,  14'd1615,  14'd654,  -14'd628,  14'd555,  14'd356,  -14'd242,  14'd1048,  14'd49,  -14'd24,  
-14'd775,  -14'd1559,  -14'd771,  -14'd594,  14'd1240,  -14'd1272,  14'd354,  -14'd844,  -14'd1877,  14'd161,  -14'd58,  -14'd72,  -14'd983,  -14'd164,  -14'd1810,  -14'd670,  
-14'd1673,  -14'd2263,  14'd618,  -14'd316,  -14'd889,  -14'd369,  -14'd572,  -14'd877,  -14'd883,  -14'd1485,  -14'd324,  -14'd743,  14'd345,  -14'd350,  -14'd1906,  -14'd506,  

-14'd12,  14'd410,  14'd649,  14'd239,  14'd363,  14'd815,  -14'd1224,  14'd983,  -14'd486,  14'd1105,  -14'd685,  -14'd722,  14'd269,  14'd304,  14'd364,  14'd304,  
14'd735,  -14'd203,  14'd18,  -14'd97,  14'd1195,  14'd928,  -14'd1213,  14'd30,  -14'd437,  -14'd606,  -14'd1188,  -14'd611,  -14'd491,  14'd719,  14'd535,  14'd306,  
14'd567,  -14'd413,  -14'd548,  14'd388,  -14'd275,  -14'd201,  14'd512,  -14'd624,  -14'd316,  -14'd824,  14'd729,  -14'd1638,  -14'd1257,  -14'd375,  14'd268,  14'd165,  
-14'd1113,  -14'd469,  -14'd167,  -14'd1356,  -14'd243,  14'd341,  -14'd307,  -14'd295,  -14'd675,  14'd704,  -14'd959,  -14'd868,  -14'd350,  14'd772,  14'd882,  -14'd1248,  
14'd682,  -14'd1602,  -14'd780,  -14'd903,  -14'd194,  14'd258,  -14'd815,  -14'd765,  14'd226,  14'd429,  14'd522,  -14'd1336,  -14'd1156,  -14'd109,  -14'd945,  14'd1289,  
-14'd865,  -14'd1233,  14'd461,  -14'd384,  -14'd706,  14'd39,  -14'd406,  14'd419,  14'd315,  14'd1119,  -14'd426,  14'd607,  14'd332,  -14'd1079,  -14'd60,  14'd102,  
14'd280,  -14'd36,  -14'd672,  -14'd1244,  -14'd1482,  14'd1364,  14'd70,  14'd97,  -14'd1019,  14'd182,  14'd68,  -14'd683,  -14'd314,  -14'd484,  -14'd937,  14'd356,  
-14'd1588,  -14'd1011,  14'd174,  -14'd1194,  -14'd180,  -14'd431,  -14'd913,  14'd574,  14'd53,  -14'd976,  -14'd403,  -14'd431,  -14'd193,  -14'd542,  14'd1403,  -14'd415,  
14'd287,  -14'd301,  -14'd448,  -14'd1047,  14'd281,  -14'd750,  -14'd1267,  -14'd973,  -14'd651,  -14'd1147,  14'd1436,  -14'd1073,  -14'd1263,  -14'd512,  -14'd806,  -14'd286,  
-14'd1197,  -14'd142,  14'd607,  -14'd710,  -14'd74,  -14'd467,  -14'd1375,  14'd1243,  -14'd809,  14'd332,  -14'd162,  -14'd1077,  -14'd1564,  -14'd330,  -14'd1302,  14'd31,  
-14'd1065,  -14'd62,  14'd127,  -14'd614,  14'd1039,  -14'd333,  -14'd614,  -14'd100,  14'd291,  -14'd1107,  14'd120,  14'd53,  -14'd1194,  14'd1338,  -14'd473,  -14'd241,  
-14'd54,  -14'd1476,  -14'd659,  -14'd1025,  14'd116,  -14'd258,  14'd344,  -14'd1167,  14'd911,  -14'd995,  -14'd625,  14'd1338,  -14'd629,  -14'd291,  -14'd75,  14'd456,  
-14'd924,  14'd1077,  -14'd20,  -14'd671,  14'd525,  14'd376,  14'd321,  14'd303,  -14'd1541,  14'd234,  -14'd416,  -14'd525,  14'd272,  -14'd580,  14'd412,  14'd460,  
-14'd204,  14'd144,  -14'd920,  -14'd1364,  14'd987,  -14'd309,  -14'd877,  -14'd457,  -14'd33,  -14'd1692,  -14'd942,  -14'd730,  -14'd936,  -14'd1071,  -14'd660,  14'd883,  
-14'd579,  14'd816,  -14'd867,  14'd1295,  14'd849,  -14'd417,  14'd587,  14'd73,  -14'd800,  -14'd561,  14'd915,  14'd195,  -14'd383,  -14'd467,  -14'd619,  14'd422,  
14'd323,  14'd37,  14'd574,  14'd229,  14'd189,  14'd887,  -14'd499,  -14'd414,  -14'd369,  -14'd1539,  -14'd413,  -14'd334,  -14'd1422,  -14'd928,  14'd354,  14'd1226,  
-14'd602,  -14'd181,  -14'd57,  -14'd1062,  14'd633,  -14'd384,  -14'd130,  14'd216,  -14'd358,  -14'd366,  14'd899,  -14'd1272,  14'd1203,  -14'd1232,  -14'd917,  14'd1407,  
14'd557,  -14'd131,  -14'd866,  14'd233,  -14'd1188,  -14'd787,  -14'd702,  14'd382,  14'd153,  -14'd8,  -14'd1388,  -14'd786,  -14'd546,  14'd412,  -14'd947,  -14'd434,  
-14'd898,  -14'd5,  -14'd1022,  14'd818,  -14'd508,  -14'd1144,  14'd641,  14'd754,  14'd414,  -14'd564,  -14'd189,  -14'd216,  14'd915,  14'd694,  -14'd1092,  -14'd832,  
-14'd684,  14'd414,  -14'd592,  -14'd642,  -14'd1197,  -14'd340,  14'd603,  -14'd1175,  -14'd181,  -14'd428,  -14'd426,  14'd435,  -14'd22,  14'd590,  14'd287,  -14'd1356,  
14'd213,  -14'd311,  -14'd662,  -14'd1246,  -14'd141,  -14'd472,  14'd1261,  14'd116,  14'd1492,  14'd236,  -14'd734,  14'd529,  -14'd602,  -14'd427,  -14'd27,  14'd255,  
-14'd13,  14'd429,  -14'd814,  -14'd541,  -14'd511,  14'd893,  14'd174,  14'd908,  14'd371,  14'd274,  14'd608,  14'd430,  14'd130,  -14'd202,  14'd346,  14'd604,  
-14'd285,  -14'd486,  -14'd414,  14'd169,  14'd33,  14'd97,  14'd120,  14'd642,  14'd203,  14'd267,  14'd813,  14'd502,  -14'd1383,  -14'd206,  14'd270,  -14'd404,  
14'd612,  -14'd891,  -14'd1310,  -14'd1674,  -14'd1126,  -14'd687,  -14'd470,  -14'd543,  -14'd650,  14'd163,  -14'd320,  -14'd1161,  14'd517,  -14'd1480,  -14'd749,  -14'd214,  
14'd1250,  14'd254,  14'd161,  -14'd333,  14'd305,  -14'd679,  -14'd727,  -14'd251,  -14'd1108,  14'd31,  14'd1107,  -14'd37,  -14'd777,  -14'd87,  -14'd1113,  14'd677,  

14'd710,  14'd297,  -14'd1423,  -14'd743,  -14'd2188,  -14'd1110,  14'd1944,  -14'd2278,  14'd57,  -14'd1118,  -14'd1470,  -14'd1409,  -14'd954,  14'd866,  -14'd1887,  -14'd1148,  
14'd944,  -14'd246,  14'd1256,  -14'd321,  -14'd284,  -14'd385,  14'd291,  14'd702,  -14'd1187,  -14'd1069,  -14'd1442,  -14'd647,  -14'd1280,  14'd1441,  14'd224,  -14'd2224,  
14'd826,  14'd914,  14'd797,  14'd925,  14'd231,  -14'd1272,  14'd553,  14'd658,  14'd354,  14'd269,  14'd1125,  14'd288,  14'd424,  -14'd1395,  -14'd882,  -14'd2041,  
14'd21,  14'd827,  14'd248,  14'd1729,  -14'd2220,  14'd489,  14'd1175,  14'd1205,  14'd588,  14'd245,  14'd1160,  14'd201,  14'd408,  14'd110,  14'd820,  -14'd1297,  
-14'd323,  14'd705,  -14'd54,  14'd2047,  -14'd247,  14'd558,  14'd280,  14'd666,  -14'd422,  -14'd386,  14'd623,  -14'd693,  14'd941,  14'd125,  -14'd197,  14'd65,  
-14'd1619,  -14'd1567,  -14'd1108,  -14'd920,  -14'd1659,  -14'd1748,  14'd447,  -14'd1806,  -14'd928,  14'd303,  14'd467,  -14'd1064,  -14'd65,  14'd451,  -14'd962,  -14'd1458,  
14'd874,  -14'd265,  14'd1296,  -14'd855,  -14'd1175,  14'd958,  -14'd62,  14'd687,  14'd19,  -14'd298,  -14'd544,  -14'd551,  14'd386,  14'd1778,  -14'd152,  -14'd155,  
-14'd896,  -14'd481,  14'd527,  -14'd247,  -14'd55,  14'd628,  14'd569,  14'd1788,  14'd1506,  14'd976,  14'd722,  -14'd212,  -14'd680,  -14'd2175,  14'd309,  -14'd507,  
-14'd620,  14'd68,  14'd359,  14'd1853,  14'd1007,  -14'd358,  14'd385,  14'd1111,  14'd962,  14'd1260,  14'd580,  -14'd1408,  14'd1675,  14'd100,  -14'd637,  14'd775,  
-14'd1656,  -14'd189,  -14'd929,  -14'd477,  -14'd16,  -14'd641,  -14'd2206,  -14'd557,  -14'd1295,  14'd776,  14'd1384,  14'd516,  14'd586,  -14'd691,  14'd576,  14'd367,  
-14'd54,  -14'd2097,  14'd1022,  -14'd460,  -14'd299,  14'd525,  -14'd1417,  14'd651,  14'd769,  -14'd959,  -14'd929,  14'd397,  -14'd761,  14'd1727,  -14'd291,  -14'd804,  
-14'd84,  -14'd1550,  14'd2413,  -14'd931,  -14'd1146,  14'd275,  14'd448,  14'd1,  -14'd1281,  -14'd164,  14'd306,  -14'd4,  14'd98,  14'd11,  14'd459,  14'd757,  
-14'd983,  -14'd322,  14'd21,  -14'd300,  -14'd542,  14'd181,  14'd288,  14'd92,  -14'd1311,  14'd678,  -14'd631,  -14'd840,  14'd887,  -14'd440,  14'd492,  -14'd117,  
-14'd2035,  -14'd1055,  14'd2051,  -14'd966,  -14'd174,  -14'd1418,  -14'd138,  -14'd133,  -14'd87,  14'd11,  14'd539,  14'd758,  -14'd1690,  14'd327,  -14'd5,  -14'd297,  
-14'd2672,  14'd1756,  14'd351,  -14'd76,  14'd53,  14'd526,  -14'd81,  -14'd32,  14'd64,  -14'd255,  14'd1157,  -14'd779,  -14'd2837,  -14'd634,  -14'd691,  -14'd1201,  
-14'd399,  14'd391,  -14'd1264,  -14'd274,  14'd1553,  14'd483,  -14'd2748,  -14'd811,  -14'd555,  14'd218,  -14'd775,  -14'd987,  -14'd680,  14'd14,  -14'd57,  -14'd1006,  
14'd155,  -14'd931,  14'd600,  14'd1033,  14'd637,  -14'd490,  -14'd705,  -14'd360,  -14'd2588,  -14'd210,  -14'd1683,  14'd559,  -14'd336,  14'd533,  14'd117,  14'd326,  
14'd875,  14'd347,  14'd904,  -14'd129,  -14'd695,  14'd189,  14'd1311,  -14'd23,  -14'd285,  -14'd908,  -14'd1161,  -14'd245,  14'd414,  14'd1442,  14'd879,  -14'd135,  
-14'd1421,  -14'd779,  14'd1637,  14'd1037,  -14'd172,  -14'd637,  14'd1209,  14'd1657,  14'd587,  -14'd856,  -14'd77,  -14'd656,  -14'd554,  -14'd744,  -14'd729,  -14'd351,  
-14'd190,  14'd506,  14'd2198,  -14'd1732,  -14'd533,  -14'd394,  -14'd791,  14'd597,  -14'd137,  -14'd1057,  -14'd363,  -14'd1286,  -14'd500,  14'd577,  -14'd1098,  -14'd1432,  
-14'd1833,  14'd219,  -14'd1256,  14'd1506,  14'd256,  14'd221,  14'd228,  14'd853,  14'd1317,  14'd244,  14'd1049,  -14'd451,  14'd377,  -14'd2054,  14'd114,  -14'd407,  
14'd452,  -14'd471,  14'd78,  14'd922,  14'd878,  -14'd308,  -14'd715,  -14'd780,  14'd1320,  14'd5,  14'd1694,  -14'd216,  14'd413,  -14'd1957,  -14'd127,  -14'd145,  
14'd977,  14'd991,  14'd1078,  -14'd25,  14'd755,  14'd183,  -14'd683,  14'd97,  -14'd584,  14'd1313,  14'd106,  14'd273,  -14'd1364,  14'd1424,  14'd435,  -14'd314,  
-14'd1599,  14'd38,  14'd225,  14'd1302,  -14'd1089,  -14'd712,  14'd1278,  -14'd242,  -14'd763,  -14'd1156,  14'd702,  -14'd716,  -14'd503,  -14'd1283,  14'd115,  -14'd476,  
-14'd972,  -14'd1861,  -14'd1674,  -14'd760,  -14'd1720,  -14'd2639,  14'd820,  -14'd1157,  14'd705,  -14'd181,  -14'd1303,  -14'd317,  -14'd648,  14'd764,  -14'd450,  -14'd1612,  

14'd78,  14'd460,  14'd1269,  14'd939,  -14'd669,  -14'd1608,  14'd630,  -14'd168,  -14'd508,  -14'd71,  14'd1057,  -14'd1186,  -14'd615,  -14'd10,  -14'd1258,  -14'd259,  
14'd704,  -14'd255,  -14'd201,  -14'd262,  -14'd1572,  14'd941,  14'd367,  -14'd718,  -14'd445,  -14'd1242,  14'd556,  -14'd814,  -14'd284,  -14'd1239,  -14'd1331,  14'd574,  
-14'd388,  14'd570,  14'd199,  14'd622,  -14'd1259,  -14'd874,  -14'd90,  -14'd855,  14'd47,  -14'd701,  14'd455,  14'd687,  -14'd221,  14'd499,  14'd313,  14'd21,  
-14'd574,  14'd808,  -14'd1040,  14'd57,  14'd921,  -14'd1765,  14'd418,  -14'd67,  -14'd677,  -14'd1131,  14'd1126,  14'd203,  14'd0,  -14'd461,  14'd623,  14'd105,  
14'd605,  14'd693,  -14'd782,  -14'd93,  14'd1061,  -14'd311,  -14'd556,  -14'd209,  14'd296,  14'd478,  14'd1216,  -14'd922,  -14'd50,  14'd859,  -14'd894,  14'd924,  
-14'd1169,  -14'd742,  14'd390,  -14'd113,  -14'd846,  -14'd639,  14'd513,  -14'd214,  -14'd272,  14'd743,  14'd596,  -14'd762,  -14'd740,  14'd479,  -14'd515,  14'd32,  
14'd555,  -14'd514,  -14'd49,  -14'd909,  -14'd870,  -14'd115,  -14'd733,  -14'd718,  -14'd375,  -14'd110,  14'd1152,  -14'd538,  -14'd850,  14'd451,  14'd138,  -14'd623,  
-14'd322,  14'd332,  -14'd627,  -14'd972,  14'd788,  -14'd336,  -14'd578,  -14'd969,  -14'd147,  14'd49,  -14'd254,  14'd604,  -14'd782,  14'd1396,  -14'd1616,  -14'd1512,  
-14'd1293,  14'd518,  -14'd1150,  14'd353,  -14'd248,  -14'd691,  -14'd752,  14'd647,  -14'd647,  -14'd1198,  -14'd1724,  -14'd125,  -14'd30,  14'd224,  -14'd26,  14'd192,  
14'd227,  14'd1104,  -14'd493,  14'd627,  -14'd1046,  -14'd347,  -14'd8,  -14'd1084,  14'd1163,  -14'd305,  14'd151,  -14'd1266,  -14'd146,  14'd307,  14'd949,  -14'd642,  
-14'd1170,  14'd312,  14'd581,  -14'd1295,  14'd147,  -14'd131,  -14'd1250,  14'd653,  -14'd252,  14'd329,  -14'd739,  -14'd564,  14'd216,  -14'd1182,  -14'd665,  -14'd16,  
-14'd926,  -14'd1614,  -14'd22,  -14'd339,  -14'd1633,  -14'd1248,  -14'd581,  -14'd1391,  -14'd622,  -14'd557,  -14'd91,  14'd785,  14'd162,  -14'd136,  -14'd311,  14'd530,  
-14'd451,  -14'd437,  14'd887,  -14'd790,  -14'd1294,  -14'd1156,  14'd387,  -14'd125,  -14'd46,  -14'd658,  -14'd976,  -14'd1611,  -14'd147,  -14'd171,  -14'd584,  -14'd309,  
14'd81,  14'd665,  -14'd994,  14'd1160,  -14'd924,  -14'd241,  -14'd1039,  -14'd580,  14'd449,  -14'd28,  -14'd388,  -14'd617,  14'd421,  14'd484,  -14'd108,  14'd688,  
-14'd436,  14'd419,  -14'd61,  -14'd450,  14'd17,  14'd117,  -14'd458,  14'd469,  -14'd976,  -14'd353,  -14'd1457,  -14'd1453,  14'd306,  14'd1021,  14'd135,  14'd431,  
-14'd422,  14'd82,  -14'd219,  14'd1070,  14'd863,  -14'd72,  -14'd357,  -14'd737,  14'd332,  -14'd652,  14'd1003,  14'd1040,  -14'd229,  -14'd415,  -14'd1003,  14'd672,  
14'd337,  -14'd36,  -14'd910,  -14'd5,  14'd55,  -14'd1288,  -14'd73,  14'd417,  14'd420,  -14'd317,  -14'd943,  -14'd636,  -14'd953,  -14'd224,  -14'd645,  14'd594,  
14'd568,  -14'd42,  -14'd912,  14'd855,  14'd210,  14'd312,  14'd180,  14'd87,  -14'd360,  14'd1188,  14'd1441,  -14'd1439,  -14'd227,  -14'd98,  -14'd940,  14'd62,  
-14'd405,  -14'd328,  -14'd357,  -14'd966,  -14'd1106,  -14'd810,  -14'd914,  -14'd160,  -14'd1205,  14'd237,  14'd698,  -14'd1632,  14'd817,  -14'd1651,  14'd221,  -14'd846,  
14'd1485,  -14'd388,  14'd476,  -14'd492,  14'd438,  -14'd1300,  -14'd1164,  -14'd1408,  -14'd495,  14'd381,  14'd763,  14'd1117,  -14'd867,  14'd33,  -14'd606,  14'd131,  
-14'd164,  14'd153,  14'd397,  -14'd169,  14'd111,  14'd1324,  -14'd283,  14'd39,  -14'd283,  -14'd1257,  14'd628,  -14'd478,  14'd163,  14'd571,  14'd204,  -14'd369,  
-14'd1360,  -14'd588,  -14'd587,  -14'd300,  14'd465,  14'd201,  -14'd8,  14'd207,  -14'd1014,  -14'd942,  14'd575,  14'd358,  14'd1121,  14'd661,  -14'd1588,  14'd507,  
-14'd470,  -14'd191,  14'd714,  -14'd1694,  -14'd1134,  -14'd1696,  -14'd82,  14'd959,  -14'd672,  -14'd927,  14'd212,  14'd265,  -14'd645,  -14'd324,  14'd1263,  14'd139,  
-14'd79,  -14'd984,  14'd1071,  -14'd214,  -14'd1217,  -14'd687,  14'd271,  14'd187,  -14'd7,  -14'd202,  -14'd1177,  -14'd603,  14'd993,  14'd223,  14'd165,  14'd508,  
-14'd351,  -14'd1029,  14'd337,  14'd712,  -14'd28,  14'd112,  -14'd51,  14'd143,  -14'd267,  -14'd436,  -14'd558,  14'd280,  14'd576,  -14'd770,  14'd516,  14'd408,  

-14'd413,  -14'd1572,  14'd141,  14'd159,  -14'd128,  -14'd646,  14'd1141,  14'd1566,  14'd826,  14'd314,  14'd592,  -14'd1692,  14'd682,  -14'd701,  14'd790,  14'd308,  
14'd1027,  14'd322,  -14'd11,  -14'd1219,  14'd1147,  -14'd91,  -14'd176,  14'd1646,  -14'd303,  14'd1194,  14'd1007,  -14'd112,  14'd1700,  -14'd1113,  14'd796,  -14'd1496,  
14'd12,  -14'd1221,  14'd251,  14'd914,  -14'd1074,  14'd560,  14'd5,  -14'd280,  14'd1,  14'd41,  -14'd265,  14'd614,  14'd1331,  -14'd808,  14'd47,  -14'd181,  
14'd1841,  -14'd50,  14'd1195,  -14'd145,  -14'd754,  -14'd1113,  14'd466,  14'd266,  14'd1320,  -14'd1186,  14'd57,  -14'd683,  14'd1961,  -14'd951,  14'd1619,  -14'd151,  
-14'd537,  -14'd911,  14'd522,  -14'd1212,  -14'd346,  -14'd839,  -14'd1060,  14'd1296,  14'd110,  -14'd201,  14'd863,  14'd825,  14'd823,  -14'd830,  -14'd739,  14'd13,  
-14'd117,  14'd824,  14'd681,  14'd1117,  14'd1494,  -14'd711,  -14'd1710,  -14'd630,  -14'd226,  -14'd152,  -14'd239,  14'd147,  -14'd191,  -14'd69,  -14'd1415,  -14'd208,  
-14'd1432,  14'd1755,  14'd129,  -14'd595,  -14'd652,  14'd1032,  -14'd1018,  -14'd1011,  14'd1103,  -14'd112,  -14'd310,  -14'd344,  14'd15,  -14'd12,  -14'd963,  -14'd815,  
-14'd1465,  14'd1644,  -14'd411,  14'd465,  14'd921,  14'd738,  14'd158,  -14'd1,  -14'd468,  14'd400,  14'd963,  -14'd403,  14'd770,  14'd379,  14'd528,  14'd1563,  
-14'd686,  14'd1457,  -14'd98,  14'd53,  14'd513,  -14'd868,  -14'd1175,  -14'd107,  14'd340,  -14'd793,  14'd578,  -14'd132,  14'd909,  14'd290,  14'd616,  14'd338,  
-14'd774,  14'd444,  14'd343,  14'd671,  -14'd996,  14'd516,  -14'd1407,  -14'd966,  -14'd229,  14'd660,  -14'd903,  14'd2147,  14'd1071,  -14'd481,  14'd604,  14'd1383,  
-14'd338,  14'd253,  14'd29,  -14'd1008,  -14'd15,  -14'd167,  -14'd1089,  14'd82,  14'd920,  -14'd1008,  14'd2262,  14'd897,  14'd329,  14'd49,  14'd777,  -14'd1059,  
14'd1087,  14'd873,  14'd1783,  -14'd1264,  -14'd498,  -14'd796,  -14'd121,  -14'd1305,  14'd795,  14'd149,  14'd141,  -14'd100,  -14'd1057,  -14'd68,  -14'd1087,  14'd862,  
14'd383,  14'd236,  -14'd537,  14'd10,  -14'd220,  -14'd455,  14'd202,  -14'd255,  -14'd678,  -14'd376,  14'd33,  -14'd1103,  14'd222,  14'd558,  14'd180,  14'd16,  
-14'd903,  14'd679,  -14'd845,  -14'd812,  14'd1908,  14'd936,  14'd113,  -14'd1089,  -14'd772,  14'd338,  14'd303,  14'd765,  14'd888,  -14'd61,  -14'd91,  14'd124,  
14'd142,  14'd488,  14'd2776,  14'd514,  14'd1642,  -14'd1708,  14'd447,  14'd96,  14'd643,  14'd1425,  14'd838,  14'd1177,  -14'd761,  14'd32,  14'd106,  14'd1364,  
14'd1294,  14'd413,  14'd407,  -14'd959,  -14'd278,  -14'd1385,  14'd697,  14'd44,  -14'd283,  -14'd932,  14'd909,  -14'd396,  -14'd1146,  14'd167,  14'd168,  14'd3,  
14'd1231,  14'd176,  14'd87,  14'd97,  14'd404,  -14'd899,  14'd938,  -14'd525,  14'd406,  14'd604,  -14'd631,  14'd471,  14'd620,  14'd1172,  -14'd728,  -14'd296,  
-14'd350,  -14'd287,  14'd528,  -14'd1309,  -14'd511,  14'd883,  14'd703,  14'd270,  14'd639,  -14'd1400,  -14'd178,  14'd1504,  14'd96,  -14'd691,  -14'd592,  -14'd886,  
-14'd201,  -14'd950,  14'd8,  -14'd243,  -14'd915,  14'd746,  14'd937,  -14'd425,  -14'd422,  -14'd454,  -14'd564,  14'd503,  14'd415,  14'd380,  -14'd1655,  14'd56,  
-14'd521,  14'd101,  14'd1490,  14'd568,  -14'd1546,  14'd343,  14'd982,  14'd829,  14'd577,  -14'd741,  -14'd381,  -14'd447,  14'd1166,  -14'd454,  14'd802,  -14'd1076,  
-14'd428,  -14'd82,  14'd362,  14'd536,  -14'd613,  -14'd307,  -14'd96,  14'd1036,  -14'd351,  -14'd138,  -14'd1048,  -14'd1213,  14'd405,  14'd1259,  -14'd427,  14'd1110,  
14'd280,  -14'd31,  14'd765,  14'd668,  -14'd850,  14'd697,  -14'd1211,  14'd1259,  -14'd1073,  14'd1161,  14'd238,  14'd801,  14'd443,  14'd496,  14'd1817,  -14'd198,  
14'd1179,  14'd317,  -14'd524,  14'd119,  14'd317,  14'd652,  -14'd622,  -14'd997,  14'd762,  -14'd604,  14'd1161,  14'd420,  14'd242,  -14'd197,  -14'd1035,  -14'd395,  
14'd236,  -14'd428,  14'd689,  -14'd1433,  14'd294,  -14'd477,  14'd1118,  -14'd683,  -14'd874,  14'd108,  -14'd63,  14'd567,  -14'd528,  14'd462,  -14'd194,  14'd529,  
14'd775,  14'd420,  14'd1611,  -14'd1174,  -14'd1195,  -14'd188,  14'd6,  -14'd219,  14'd174,  -14'd203,  -14'd1002,  -14'd562,  -14'd1737,  14'd1321,  -14'd818,  -14'd579,  

14'd204,  14'd1036,  14'd529,  -14'd247,  14'd380,  14'd274,  14'd1077,  14'd527,  -14'd354,  -14'd49,  14'd405,  -14'd6,  14'd629,  14'd665,  14'd1409,  -14'd13,  
14'd2099,  14'd435,  14'd1675,  -14'd453,  -14'd968,  14'd475,  14'd1491,  -14'd757,  -14'd28,  -14'd1232,  14'd1007,  14'd739,  -14'd82,  14'd1588,  -14'd468,  14'd1147,  
14'd578,  -14'd429,  14'd1390,  -14'd795,  -14'd1148,  -14'd869,  14'd2068,  -14'd1479,  -14'd1705,  -14'd858,  14'd619,  -14'd1497,  14'd261,  14'd320,  -14'd1445,  -14'd712,  
-14'd777,  -14'd45,  -14'd2689,  -14'd2054,  -14'd164,  -14'd1356,  14'd1892,  -14'd1467,  -14'd1048,  -14'd2254,  14'd1773,  -14'd45,  -14'd322,  14'd1174,  -14'd836,  -14'd172,  
-14'd979,  14'd290,  -14'd2203,  -14'd1186,  -14'd1358,  -14'd881,  -14'd2274,  -14'd2198,  -14'd1974,  -14'd557,  -14'd120,  -14'd1408,  -14'd2081,  -14'd323,  -14'd1100,  14'd934,  
14'd1708,  -14'd123,  14'd579,  -14'd12,  -14'd818,  -14'd954,  14'd59,  14'd67,  14'd1447,  -14'd1200,  14'd1365,  14'd1306,  14'd1994,  14'd104,  14'd889,  14'd258,  
-14'd63,  14'd1136,  -14'd443,  -14'd1205,  14'd830,  -14'd1106,  14'd847,  14'd18,  -14'd1040,  14'd1222,  14'd955,  -14'd604,  -14'd140,  14'd547,  14'd158,  14'd147,  
-14'd312,  -14'd1596,  14'd578,  -14'd610,  -14'd619,  -14'd2931,  -14'd198,  -14'd1152,  14'd351,  -14'd72,  14'd221,  14'd708,  -14'd357,  -14'd1047,  -14'd1418,  -14'd1419,  
14'd349,  14'd337,  -14'd1133,  -14'd184,  -14'd1128,  14'd253,  -14'd629,  -14'd2188,  14'd1655,  14'd1427,  -14'd779,  -14'd949,  -14'd604,  -14'd722,  -14'd1236,  -14'd1366,  
14'd1673,  -14'd1808,  -14'd24,  14'd1004,  14'd1254,  -14'd426,  -14'd12,  -14'd1804,  14'd476,  14'd1372,  -14'd1349,  14'd1770,  14'd181,  14'd68,  -14'd793,  14'd157,  
-14'd766,  14'd55,  14'd1345,  14'd279,  -14'd900,  -14'd1001,  14'd748,  -14'd223,  -14'd462,  14'd70,  -14'd8,  -14'd596,  -14'd1296,  14'd21,  -14'd1071,  14'd657,  
-14'd1227,  14'd1433,  14'd1752,  -14'd1219,  -14'd579,  -14'd759,  14'd270,  -14'd296,  14'd448,  -14'd694,  -14'd948,  -14'd1451,  -14'd1415,  14'd1254,  14'd251,  -14'd2178,  
14'd951,  -14'd2397,  14'd846,  14'd184,  -14'd1334,  -14'd914,  -14'd1378,  -14'd962,  -14'd1063,  14'd386,  -14'd979,  -14'd106,  -14'd2435,  -14'd64,  -14'd595,  14'd363,  
14'd1650,  -14'd566,  -14'd2114,  14'd536,  14'd72,  14'd977,  -14'd979,  -14'd205,  14'd1777,  14'd306,  14'd1827,  14'd844,  14'd733,  -14'd39,  -14'd255,  14'd1114,  
14'd1121,  14'd638,  14'd312,  14'd509,  14'd1400,  14'd1305,  14'd946,  -14'd221,  14'd1034,  14'd1015,  14'd2212,  14'd1156,  14'd748,  -14'd205,  14'd957,  14'd687,  
-14'd828,  14'd433,  -14'd1172,  -14'd9,  14'd1008,  -14'd619,  14'd361,  14'd595,  14'd693,  -14'd1680,  -14'd733,  -14'd827,  14'd848,  -14'd374,  14'd454,  14'd530,  
14'd116,  -14'd762,  14'd635,  14'd528,  -14'd617,  14'd1111,  -14'd513,  14'd657,  -14'd634,  -14'd210,  14'd846,  -14'd255,  14'd131,  14'd1299,  14'd53,  -14'd761,  
14'd549,  -14'd1527,  14'd1208,  14'd1068,  -14'd320,  -14'd360,  -14'd438,  14'd1036,  -14'd2131,  14'd363,  14'd929,  -14'd170,  14'd1611,  -14'd562,  14'd785,  -14'd2034,  
-14'd72,  -14'd563,  -14'd1011,  14'd1537,  14'd1467,  -14'd30,  14'd1103,  14'd940,  -14'd1721,  -14'd601,  14'd1231,  14'd818,  14'd716,  -14'd836,  14'd1478,  -14'd54,  
-14'd222,  14'd137,  -14'd540,  14'd820,  -14'd509,  14'd199,  14'd707,  14'd1753,  -14'd746,  14'd1236,  14'd766,  14'd297,  14'd1808,  -14'd272,  14'd225,  14'd777,  
14'd196,  -14'd198,  14'd151,  14'd48,  14'd935,  -14'd657,  -14'd1875,  14'd526,  14'd283,  14'd196,  14'd66,  -14'd2063,  14'd491,  -14'd100,  -14'd1348,  -14'd561,  
-14'd1730,  14'd814,  -14'd586,  14'd732,  -14'd529,  -14'd115,  -14'd2769,  14'd509,  14'd1500,  14'd333,  14'd632,  -14'd2365,  14'd1021,  14'd916,  -14'd1048,  14'd483,  
14'd38,  -14'd709,  -14'd2412,  14'd191,  -14'd917,  14'd973,  -14'd445,  14'd284,  -14'd2044,  -14'd453,  14'd1310,  14'd20,  14'd1202,  -14'd3610,  -14'd1095,  -14'd842,  
-14'd1677,  -14'd1524,  -14'd4021,  14'd131,  14'd806,  -14'd386,  -14'd466,  -14'd110,  14'd580,  -14'd1872,  14'd988,  14'd30,  14'd139,  -14'd169,  -14'd1593,  14'd4,  
14'd154,  -14'd1667,  -14'd1355,  -14'd1457,  14'd349,  -14'd2114,  -14'd1379,  14'd937,  -14'd297,  14'd2034,  14'd36,  -14'd1272,  -14'd1207,  -14'd947,  -14'd908,  14'd739,  

-14'd676,  -14'd586,  14'd1317,  14'd908,  -14'd248,  -14'd516,  -14'd1183,  14'd367,  14'd278,  -14'd394,  -14'd606,  -14'd486,  -14'd658,  -14'd633,  14'd649,  -14'd346,  
14'd1516,  -14'd925,  14'd628,  14'd1615,  14'd449,  14'd1717,  -14'd331,  14'd479,  -14'd890,  -14'd943,  -14'd1194,  14'd118,  14'd1426,  14'd586,  14'd1008,  -14'd2179,  
-14'd661,  14'd399,  -14'd368,  -14'd547,  -14'd450,  14'd1838,  -14'd640,  14'd1214,  14'd2385,  14'd1181,  -14'd65,  -14'd1221,  14'd1084,  -14'd1024,  14'd1660,  -14'd1155,  
-14'd158,  -14'd464,  -14'd954,  14'd226,  -14'd841,  -14'd836,  -14'd2012,  -14'd60,  -14'd1726,  14'd750,  -14'd967,  -14'd1297,  14'd4,  -14'd1375,  14'd487,  14'd1575,  
-14'd120,  -14'd798,  14'd711,  14'd170,  14'd561,  -14'd191,  14'd589,  14'd1260,  -14'd94,  14'd564,  -14'd85,  14'd500,  14'd53,  -14'd812,  -14'd219,  -14'd1308,  
14'd985,  -14'd161,  14'd239,  -14'd767,  -14'd1195,  14'd368,  14'd160,  -14'd512,  -14'd432,  14'd186,  -14'd130,  14'd797,  -14'd441,  14'd1290,  14'd976,  -14'd797,  
14'd637,  -14'd1064,  14'd2740,  14'd559,  -14'd155,  14'd1456,  -14'd736,  14'd257,  14'd1007,  -14'd1537,  -14'd1340,  -14'd1317,  -14'd253,  14'd75,  -14'd1359,  -14'd834,  
-14'd829,  14'd2021,  -14'd1417,  -14'd844,  14'd521,  14'd2323,  -14'd385,  14'd1560,  14'd1741,  -14'd601,  -14'd21,  14'd208,  14'd626,  14'd686,  14'd85,  14'd550,  
14'd502,  14'd650,  -14'd393,  14'd305,  14'd284,  14'd545,  -14'd1199,  14'd1095,  -14'd1156,  -14'd111,  -14'd509,  -14'd1207,  14'd882,  14'd498,  14'd1442,  -14'd719,  
-14'd175,  -14'd876,  14'd144,  14'd307,  14'd1303,  14'd267,  14'd48,  14'd418,  -14'd908,  14'd743,  14'd1446,  14'd2314,  14'd230,  -14'd1179,  14'd205,  14'd977,  
14'd778,  -14'd584,  14'd1439,  14'd944,  14'd231,  14'd1455,  -14'd97,  14'd268,  -14'd458,  -14'd344,  -14'd70,  14'd740,  -14'd1119,  14'd234,  -14'd889,  -14'd910,  
14'd759,  14'd1982,  -14'd45,  -14'd491,  14'd576,  14'd921,  14'd1047,  -14'd882,  -14'd8,  -14'd1236,  14'd181,  14'd326,  14'd1041,  -14'd870,  -14'd1028,  -14'd265,  
14'd538,  14'd1544,  -14'd1502,  14'd235,  14'd1282,  -14'd103,  14'd990,  -14'd1263,  -14'd870,  -14'd281,  -14'd1342,  -14'd2015,  -14'd1078,  14'd798,  14'd198,  -14'd1092,  
14'd835,  14'd1795,  -14'd893,  -14'd1897,  14'd934,  14'd14,  -14'd755,  14'd57,  -14'd407,  -14'd896,  -14'd836,  14'd221,  -14'd212,  14'd552,  14'd1507,  14'd542,  
14'd423,  14'd1269,  14'd267,  -14'd159,  14'd1151,  -14'd352,  -14'd70,  -14'd355,  -14'd739,  -14'd3395,  14'd773,  -14'd704,  14'd9,  -14'd960,  14'd547,  14'd57,  
14'd770,  -14'd583,  14'd512,  14'd1240,  14'd144,  -14'd391,  14'd201,  14'd1153,  -14'd971,  -14'd560,  -14'd1105,  -14'd131,  -14'd1016,  -14'd422,  14'd657,  -14'd254,  
14'd36,  -14'd422,  -14'd372,  -14'd1146,  -14'd346,  -14'd502,  14'd2346,  14'd1187,  -14'd196,  -14'd1666,  -14'd847,  -14'd468,  -14'd1693,  14'd190,  14'd988,  -14'd1617,  
14'd1007,  14'd629,  14'd844,  14'd489,  -14'd284,  -14'd624,  -14'd325,  -14'd238,  14'd885,  14'd100,  -14'd48,  -14'd156,  -14'd889,  14'd1481,  -14'd130,  -14'd1238,  
14'd1086,  14'd1082,  14'd383,  -14'd405,  14'd49,  14'd986,  14'd706,  -14'd208,  14'd20,  14'd524,  14'd434,  14'd1071,  14'd540,  14'd1433,  -14'd1352,  -14'd559,  
14'd827,  14'd795,  14'd1069,  -14'd663,  14'd301,  14'd1048,  14'd1034,  14'd855,  -14'd318,  -14'd436,  14'd230,  14'd447,  -14'd154,  -14'd172,  -14'd2019,  14'd512,  
-14'd1038,  14'd1060,  14'd250,  14'd3,  -14'd1405,  14'd578,  -14'd373,  14'd1138,  14'd221,  -14'd235,  -14'd286,  14'd1136,  -14'd835,  -14'd734,  -14'd855,  14'd196,  
14'd330,  -14'd319,  -14'd758,  -14'd279,  14'd137,  14'd905,  14'd262,  14'd138,  14'd265,  14'd424,  14'd14,  14'd437,  14'd817,  -14'd601,  14'd220,  -14'd279,  
-14'd597,  -14'd1484,  -14'd708,  -14'd423,  14'd399,  14'd229,  -14'd569,  -14'd205,  14'd476,  14'd180,  -14'd521,  14'd871,  -14'd103,  -14'd605,  -14'd1290,  14'd217,  
14'd2479,  -14'd1481,  14'd1738,  -14'd440,  14'd879,  14'd33,  -14'd740,  14'd516,  14'd706,  14'd544,  14'd939,  14'd1163,  14'd431,  -14'd455,  -14'd2363,  -14'd936,  
14'd2009,  14'd975,  -14'd435,  -14'd1934,  -14'd439,  -14'd1379,  -14'd989,  14'd185,  -14'd1081,  -14'd1636,  -14'd1755,  -14'd880,  14'd253,  -14'd662,  -14'd2239,  14'd514,  

14'd1503,  14'd612,  -14'd1190,  -14'd50,  -14'd451,  -14'd672,  14'd911,  -14'd682,  14'd1180,  -14'd623,  -14'd711,  14'd328,  -14'd2050,  -14'd594,  14'd547,  -14'd1354,  
14'd1045,  14'd601,  14'd191,  -14'd703,  -14'd862,  14'd15,  -14'd342,  14'd900,  -14'd501,  14'd1255,  -14'd482,  -14'd683,  -14'd227,  -14'd229,  14'd275,  -14'd352,  
14'd767,  -14'd607,  -14'd360,  14'd91,  14'd31,  14'd225,  -14'd1543,  -14'd1058,  14'd5,  14'd1703,  -14'd136,  14'd86,  -14'd1134,  -14'd412,  14'd404,  14'd1386,  
-14'd458,  -14'd910,  14'd571,  14'd693,  -14'd568,  -14'd906,  -14'd385,  -14'd657,  14'd567,  14'd302,  14'd1030,  -14'd1712,  14'd1098,  -14'd1262,  -14'd247,  14'd96,  
14'd1212,  -14'd785,  14'd218,  -14'd57,  14'd1595,  -14'd548,  -14'd648,  14'd815,  -14'd874,  -14'd655,  14'd474,  14'd378,  -14'd584,  14'd168,  -14'd37,  14'd2298,  
14'd237,  -14'd288,  14'd1078,  -14'd326,  14'd1293,  14'd629,  -14'd1016,  -14'd82,  14'd845,  14'd1655,  -14'd936,  -14'd80,  -14'd447,  -14'd738,  14'd1963,  14'd223,  
-14'd610,  14'd990,  14'd639,  14'd72,  14'd445,  -14'd497,  -14'd283,  14'd1662,  14'd214,  14'd745,  -14'd1656,  -14'd944,  14'd425,  14'd681,  14'd1563,  14'd2097,  
-14'd426,  -14'd24,  14'd230,  14'd1115,  -14'd1466,  -14'd155,  -14'd712,  14'd536,  14'd286,  -14'd943,  14'd349,  -14'd58,  14'd911,  -14'd1184,  -14'd675,  14'd113,  
-14'd996,  -14'd708,  -14'd994,  -14'd53,  -14'd824,  -14'd329,  14'd193,  14'd245,  -14'd291,  14'd246,  -14'd637,  14'd1121,  -14'd600,  -14'd1958,  -14'd710,  14'd546,  
-14'd33,  14'd1513,  -14'd881,  -14'd504,  -14'd1,  14'd754,  -14'd67,  14'd1565,  -14'd582,  14'd720,  -14'd617,  14'd668,  14'd1816,  14'd88,  -14'd1101,  14'd18,  
-14'd535,  -14'd736,  -14'd853,  14'd1693,  14'd1853,  14'd357,  -14'd3714,  14'd1268,  -14'd5,  14'd1822,  14'd67,  14'd1950,  -14'd389,  -14'd590,  -14'd126,  14'd94,  
-14'd423,  14'd2471,  14'd949,  14'd247,  -14'd59,  14'd1044,  -14'd812,  14'd200,  -14'd298,  14'd1564,  14'd1764,  14'd1037,  -14'd26,  14'd226,  -14'd138,  14'd1148,  
14'd438,  14'd61,  -14'd7,  14'd849,  -14'd748,  14'd10,  -14'd1271,  -14'd577,  -14'd187,  14'd314,  14'd1040,  14'd1412,  14'd26,  -14'd1057,  -14'd292,  14'd370,  
-14'd1172,  -14'd887,  14'd65,  -14'd844,  14'd1311,  -14'd1632,  14'd771,  14'd394,  -14'd581,  -14'd114,  14'd744,  14'd357,  14'd944,  14'd750,  -14'd100,  14'd1537,  
14'd1564,  -14'd553,  -14'd1412,  -14'd162,  14'd282,  14'd16,  -14'd551,  -14'd1421,  -14'd618,  -14'd22,  -14'd137,  -14'd591,  14'd522,  -14'd353,  -14'd429,  14'd807,  
-14'd141,  -14'd1299,  -14'd296,  14'd825,  14'd2747,  -14'd102,  -14'd1404,  14'd502,  14'd584,  14'd938,  -14'd441,  14'd1672,  -14'd348,  14'd847,  14'd982,  14'd140,  
14'd984,  14'd541,  -14'd426,  14'd700,  14'd1362,  -14'd33,  14'd271,  -14'd1705,  14'd1723,  14'd1962,  -14'd745,  14'd938,  14'd1425,  -14'd96,  -14'd265,  14'd574,  
-14'd435,  14'd1432,  14'd140,  -14'd530,  14'd335,  -14'd1645,  14'd691,  -14'd272,  14'd1448,  -14'd672,  -14'd739,  14'd515,  -14'd1250,  14'd744,  -14'd645,  -14'd1112,  
14'd439,  -14'd166,  14'd145,  -14'd1475,  14'd21,  -14'd20,  -14'd1139,  -14'd605,  -14'd183,  -14'd345,  -14'd2145,  14'd247,  14'd361,  14'd173,  -14'd633,  -14'd1573,  
-14'd700,  -14'd156,  14'd1757,  -14'd45,  -14'd308,  14'd268,  14'd282,  -14'd337,  14'd407,  14'd150,  -14'd1619,  14'd854,  -14'd656,  14'd47,  14'd787,  -14'd1598,  
14'd501,  14'd337,  -14'd25,  -14'd156,  14'd269,  14'd1541,  14'd1187,  14'd1975,  14'd675,  -14'd101,  -14'd107,  14'd1261,  14'd227,  14'd248,  14'd65,  14'd949,  
-14'd144,  -14'd233,  -14'd1092,  14'd553,  -14'd60,  -14'd149,  -14'd2002,  14'd1244,  -14'd1209,  -14'd16,  -14'd206,  -14'd1048,  14'd602,  14'd703,  14'd1047,  -14'd320,  
14'd866,  -14'd1552,  -14'd612,  -14'd384,  -14'd1152,  -14'd776,  14'd612,  -14'd328,  14'd230,  14'd1574,  14'd115,  14'd1859,  14'd433,  -14'd58,  14'd560,  -14'd742,  
14'd185,  -14'd495,  -14'd393,  14'd1169,  -14'd707,  14'd1438,  -14'd1256,  -14'd1318,  14'd523,  -14'd58,  14'd1116,  14'd1259,  -14'd2,  14'd602,  14'd211,  -14'd367,  
14'd1577,  -14'd528,  14'd2695,  14'd1303,  -14'd629,  14'd1992,  -14'd168,  14'd579,  14'd1597,  -14'd477,  -14'd231,  14'd532,  -14'd238,  14'd14,  14'd1652,  -14'd964,  

-14'd523,  14'd733,  -14'd503,  -14'd696,  -14'd204,  14'd385,  14'd389,  14'd1188,  14'd941,  -14'd138,  14'd57,  -14'd263,  14'd2208,  14'd799,  14'd190,  -14'd349,  
14'd902,  14'd1179,  14'd1827,  -14'd71,  14'd129,  14'd471,  14'd498,  14'd215,  14'd487,  14'd40,  14'd520,  -14'd1229,  14'd700,  14'd355,  14'd511,  14'd863,  
-14'd629,  -14'd726,  14'd415,  14'd643,  -14'd130,  14'd144,  14'd628,  14'd891,  14'd263,  14'd69,  -14'd305,  14'd371,  14'd522,  -14'd415,  -14'd572,  14'd966,  
14'd768,  14'd187,  14'd1264,  14'd487,  -14'd1044,  14'd599,  -14'd927,  -14'd88,  -14'd480,  -14'd337,  -14'd717,  14'd468,  14'd979,  -14'd702,  -14'd157,  14'd122,  
14'd423,  14'd790,  14'd281,  -14'd392,  -14'd556,  -14'd76,  14'd245,  -14'd18,  -14'd319,  -14'd844,  -14'd802,  14'd1000,  -14'd426,  -14'd670,  14'd553,  -14'd1254,  
-14'd948,  14'd388,  -14'd672,  14'd551,  14'd76,  14'd298,  -14'd756,  -14'd1440,  -14'd359,  -14'd1495,  14'd1026,  14'd664,  14'd15,  14'd1259,  -14'd2,  14'd930,  
-14'd434,  14'd17,  14'd1782,  -14'd818,  -14'd740,  14'd1383,  14'd1021,  -14'd1874,  -14'd16,  -14'd587,  14'd1466,  14'd115,  14'd159,  14'd693,  -14'd1233,  14'd338,  
14'd47,  14'd2255,  -14'd1128,  14'd836,  14'd542,  14'd1532,  14'd2220,  -14'd944,  14'd175,  14'd338,  14'd133,  -14'd102,  -14'd360,  14'd866,  -14'd260,  14'd1573,  
14'd5,  14'd1379,  14'd215,  -14'd1098,  14'd1780,  -14'd400,  -14'd602,  14'd524,  -14'd878,  14'd919,  -14'd114,  14'd111,  14'd1249,  -14'd677,  14'd425,  14'd197,  
14'd2388,  14'd499,  -14'd636,  -14'd1566,  -14'd604,  -14'd851,  -14'd155,  -14'd801,  14'd1297,  14'd1861,  14'd264,  14'd996,  -14'd332,  -14'd1040,  14'd459,  14'd63,  
-14'd351,  -14'd712,  -14'd331,  -14'd776,  -14'd1561,  -14'd888,  14'd787,  14'd919,  -14'd605,  -14'd163,  14'd573,  14'd681,  14'd744,  -14'd480,  14'd175,  -14'd315,  
14'd1215,  14'd450,  14'd76,  -14'd743,  14'd66,  -14'd1073,  14'd746,  -14'd689,  -14'd1097,  -14'd1126,  -14'd450,  -14'd493,  14'd49,  14'd147,  14'd256,  -14'd74,  
-14'd32,  14'd2373,  14'd658,  -14'd1385,  14'd597,  -14'd1284,  14'd1149,  -14'd83,  -14'd273,  14'd749,  -14'd1572,  -14'd407,  -14'd2503,  14'd2437,  -14'd15,  14'd1025,  
-14'd592,  14'd1181,  14'd983,  -14'd370,  14'd107,  -14'd395,  14'd370,  14'd832,  14'd76,  -14'd1134,  14'd143,  14'd116,  -14'd2210,  14'd953,  14'd279,  -14'd1471,  
14'd165,  14'd172,  14'd1013,  -14'd1751,  -14'd1573,  -14'd86,  14'd1027,  -14'd51,  -14'd350,  -14'd1013,  -14'd900,  -14'd433,  -14'd926,  -14'd927,  14'd2060,  -14'd1485,  
14'd2275,  14'd178,  14'd248,  -14'd2362,  -14'd1032,  -14'd775,  14'd77,  -14'd1451,  -14'd948,  14'd55,  -14'd1568,  14'd1082,  -14'd2663,  14'd571,  -14'd808,  14'd664,  
-14'd504,  14'd1041,  14'd868,  -14'd1102,  -14'd1472,  -14'd441,  14'd1099,  -14'd186,  14'd2557,  14'd986,  -14'd167,  14'd683,  -14'd1019,  14'd2,  14'd168,  -14'd1196,  
-14'd17,  -14'd562,  -14'd18,  -14'd131,  -14'd358,  14'd476,  -14'd395,  -14'd987,  14'd1139,  14'd1354,  -14'd1350,  -14'd839,  -14'd799,  14'd1524,  -14'd633,  -14'd2387,  
-14'd292,  -14'd200,  -14'd1308,  14'd240,  -14'd103,  -14'd634,  -14'd549,  -14'd99,  14'd988,  14'd619,  -14'd1702,  14'd260,  -14'd739,  -14'd16,  -14'd829,  -14'd360,  
14'd457,  -14'd18,  -14'd479,  14'd480,  -14'd109,  14'd1185,  -14'd1704,  -14'd104,  14'd685,  -14'd213,  -14'd466,  -14'd1286,  -14'd684,  -14'd626,  -14'd319,  -14'd1252,  
14'd1977,  -14'd563,  14'd721,  -14'd110,  -14'd3726,  14'd1409,  -14'd961,  -14'd170,  14'd327,  -14'd715,  -14'd785,  14'd2428,  -14'd166,  14'd1802,  14'd1130,  -14'd711,  
14'd619,  -14'd387,  14'd1050,  -14'd153,  -14'd135,  14'd897,  14'd2344,  14'd876,  -14'd96,  14'd863,  14'd345,  14'd381,  14'd290,  14'd1241,  14'd1163,  -14'd423,  
14'd29,  -14'd995,  -14'd526,  -14'd482,  14'd610,  -14'd672,  14'd352,  14'd821,  14'd830,  -14'd1475,  14'd456,  -14'd1399,  -14'd537,  14'd89,  -14'd247,  14'd164,  
-14'd43,  -14'd544,  14'd767,  14'd1054,  -14'd612,  -14'd885,  14'd293,  14'd124,  -14'd393,  -14'd557,  14'd132,  -14'd1466,  14'd653,  -14'd153,  -14'd1148,  -14'd422,  
-14'd1483,  -14'd1401,  -14'd961,  -14'd116,  14'd449,  -14'd888,  14'd162,  -14'd305,  14'd398,  14'd1697,  -14'd994,  -14'd225,  14'd1278,  -14'd797,  -14'd1087,  14'd858,  

14'd806,  14'd1088,  -14'd1176,  -14'd985,  14'd1272,  -14'd1033,  -14'd1251,  14'd1783,  -14'd658,  14'd593,  14'd23,  14'd175,  14'd1236,  14'd134,  -14'd1305,  14'd1207,  
-14'd630,  -14'd726,  -14'd953,  14'd652,  14'd1213,  -14'd723,  -14'd2051,  14'd1334,  14'd231,  14'd147,  -14'd132,  14'd620,  14'd347,  14'd715,  14'd1072,  14'd212,  
14'd1178,  -14'd628,  -14'd306,  -14'd209,  -14'd1240,  14'd1130,  14'd643,  -14'd1379,  14'd227,  -14'd1271,  14'd2313,  14'd129,  14'd655,  14'd719,  -14'd145,  14'd1134,  
-14'd870,  -14'd732,  -14'd650,  14'd339,  -14'd215,  14'd26,  14'd2047,  -14'd860,  -14'd862,  14'd239,  14'd407,  14'd365,  14'd1010,  -14'd856,  14'd698,  -14'd472,  
-14'd356,  14'd159,  14'd64,  -14'd989,  -14'd1133,  -14'd617,  14'd1036,  14'd265,  -14'd680,  -14'd1643,  14'd221,  -14'd913,  -14'd1134,  14'd1727,  14'd714,  14'd14,  
14'd31,  14'd157,  -14'd1532,  -14'd116,  14'd233,  -14'd1558,  -14'd1754,  -14'd244,  -14'd620,  14'd528,  14'd1666,  -14'd237,  -14'd293,  14'd172,  14'd149,  -14'd544,  
14'd1260,  -14'd241,  14'd1170,  14'd195,  14'd230,  -14'd885,  -14'd81,  -14'd1422,  -14'd1462,  14'd891,  14'd1047,  14'd1707,  14'd429,  -14'd441,  14'd617,  14'd689,  
-14'd544,  -14'd677,  14'd395,  14'd219,  14'd1025,  -14'd1918,  -14'd880,  14'd267,  -14'd999,  14'd1934,  14'd1902,  14'd1088,  -14'd160,  -14'd6,  14'd877,  -14'd204,  
-14'd404,  -14'd76,  -14'd671,  -14'd1171,  -14'd817,  -14'd2168,  14'd516,  -14'd491,  -14'd927,  14'd1495,  14'd34,  -14'd528,  14'd1441,  -14'd38,  -14'd711,  14'd393,  
-14'd917,  14'd1304,  14'd1192,  -14'd1463,  14'd290,  -14'd111,  -14'd214,  14'd1608,  -14'd1721,  14'd2112,  -14'd644,  14'd1054,  -14'd1375,  14'd335,  -14'd1738,  -14'd754,  
-14'd1458,  -14'd1352,  -14'd708,  -14'd1289,  -14'd442,  14'd211,  -14'd1013,  -14'd1320,  14'd987,  14'd1178,  14'd604,  -14'd169,  14'd297,  14'd579,  -14'd411,  14'd729,  
14'd197,  -14'd1410,  -14'd376,  14'd1062,  14'd248,  -14'd647,  -14'd2063,  -14'd273,  14'd472,  14'd661,  -14'd444,  14'd106,  -14'd744,  14'd326,  -14'd1424,  14'd1206,  
14'd690,  -14'd1607,  14'd195,  14'd1033,  14'd444,  -14'd58,  14'd87,  14'd227,  14'd1454,  14'd1855,  -14'd1030,  14'd513,  -14'd809,  -14'd1232,  -14'd999,  14'd635,  
-14'd2120,  14'd293,  -14'd392,  -14'd33,  14'd1391,  -14'd317,  -14'd1573,  14'd506,  14'd227,  14'd1167,  -14'd951,  -14'd1216,  14'd1099,  -14'd404,  14'd1227,  14'd1250,  
-14'd662,  -14'd717,  -14'd1488,  -14'd60,  14'd738,  14'd328,  -14'd206,  -14'd965,  14'd516,  14'd1844,  -14'd147,  14'd1299,  -14'd1038,  14'd1583,  14'd138,  -14'd1278,  
-14'd790,  -14'd1714,  14'd469,  -14'd406,  14'd689,  14'd76,  -14'd1024,  -14'd845,  14'd1808,  -14'd1109,  14'd321,  -14'd1112,  14'd937,  -14'd1543,  14'd841,  14'd671,  
-14'd961,  -14'd1155,  -14'd1238,  -14'd296,  -14'd832,  14'd1575,  -14'd1559,  14'd822,  -14'd240,  14'd911,  14'd236,  14'd1611,  14'd329,  -14'd1020,  14'd347,  14'd214,  
14'd947,  -14'd630,  -14'd464,  14'd391,  -14'd796,  14'd1400,  14'd451,  14'd1274,  -14'd906,  -14'd1054,  14'd1334,  14'd992,  14'd20,  -14'd477,  -14'd27,  14'd70,  
-14'd14,  14'd1603,  -14'd320,  14'd0,  14'd737,  -14'd61,  14'd231,  14'd1301,  -14'd332,  14'd732,  -14'd232,  -14'd200,  -14'd402,  -14'd103,  -14'd179,  14'd227,  
-14'd82,  -14'd230,  14'd556,  -14'd55,  14'd1648,  14'd214,  14'd206,  14'd1750,  14'd1162,  -14'd74,  14'd72,  -14'd1500,  14'd309,  -14'd963,  14'd483,  14'd63,  
-14'd1,  -14'd571,  14'd801,  14'd1105,  14'd362,  -14'd966,  14'd749,  -14'd375,  14'd620,  14'd391,  -14'd456,  14'd649,  14'd1746,  14'd305,  14'd760,  14'd978,  
-14'd22,  -14'd408,  14'd48,  -14'd61,  -14'd1311,  -14'd603,  14'd1253,  14'd365,  14'd845,  -14'd1852,  14'd577,  14'd433,  14'd1063,  -14'd1365,  14'd1380,  14'd877,  
14'd1457,  -14'd229,  -14'd1175,  14'd542,  14'd615,  14'd383,  -14'd1479,  -14'd85,  -14'd1122,  14'd849,  14'd1348,  14'd256,  14'd1428,  -14'd922,  -14'd488,  -14'd862,  
14'd504,  14'd2175,  -14'd497,  14'd1160,  -14'd49,  -14'd484,  -14'd573,  14'd417,  14'd144,  -14'd98,  -14'd190,  14'd1402,  14'd490,  -14'd1012,  14'd7,  -14'd601,  
14'd2026,  14'd1455,  14'd799,  -14'd443,  -14'd130,  14'd572,  14'd356,  14'd186,  14'd1995,  14'd3185,  -14'd1120,  14'd2041,  14'd1153,  14'd1414,  14'd1028,  14'd828,  

14'd1337,  -14'd385,  -14'd1714,  -14'd1030,  14'd699,  -14'd124,  14'd714,  14'd544,  -14'd504,  14'd494,  14'd286,  -14'd628,  -14'd2184,  14'd530,  14'd928,  -14'd457,  
-14'd1170,  14'd40,  -14'd2865,  14'd331,  14'd436,  14'd810,  14'd129,  -14'd153,  14'd893,  14'd213,  -14'd547,  14'd26,  -14'd1497,  -14'd1143,  -14'd707,  14'd445,  
-14'd116,  14'd308,  -14'd1192,  14'd1591,  -14'd579,  14'd1642,  -14'd276,  -14'd161,  -14'd608,  14'd1703,  14'd69,  14'd23,  14'd196,  -14'd1913,  14'd984,  14'd177,  
-14'd928,  -14'd709,  -14'd649,  14'd837,  14'd214,  14'd124,  14'd99,  -14'd433,  14'd1039,  14'd1142,  -14'd453,  -14'd441,  14'd828,  -14'd1017,  14'd214,  14'd1213,  
-14'd692,  -14'd2169,  -14'd547,  14'd853,  14'd777,  14'd256,  -14'd186,  14'd309,  -14'd163,  14'd1026,  14'd260,  -14'd487,  -14'd1747,  14'd731,  -14'd23,  14'd520,  
14'd875,  14'd615,  -14'd604,  -14'd567,  14'd73,  14'd266,  -14'd434,  14'd876,  14'd895,  14'd15,  14'd58,  14'd179,  14'd148,  14'd75,  14'd221,  14'd970,  
14'd1316,  14'd1244,  -14'd105,  -14'd1251,  -14'd676,  -14'd14,  -14'd1360,  -14'd73,  14'd982,  14'd585,  -14'd2414,  -14'd675,  14'd312,  -14'd250,  14'd160,  14'd1538,  
-14'd80,  -14'd344,  -14'd496,  -14'd587,  14'd599,  -14'd1,  14'd634,  -14'd469,  -14'd163,  14'd949,  14'd445,  14'd1908,  -14'd276,  -14'd190,  14'd1167,  14'd997,  
14'd525,  -14'd224,  -14'd2788,  14'd1249,  -14'd97,  14'd943,  -14'd439,  -14'd853,  14'd777,  14'd123,  -14'd876,  -14'd443,  -14'd234,  -14'd552,  14'd920,  14'd1179,  
-14'd1747,  -14'd1494,  -14'd1226,  14'd1581,  -14'd1617,  14'd62,  -14'd269,  14'd215,  14'd172,  -14'd2359,  14'd566,  -14'd545,  14'd1474,  14'd792,  -14'd391,  -14'd808,  
14'd175,  -14'd1009,  14'd570,  14'd456,  14'd39,  -14'd844,  -14'd1020,  14'd790,  14'd1215,  14'd396,  -14'd2017,  14'd691,  14'd1836,  -14'd306,  14'd1130,  14'd668,  
-14'd149,  -14'd561,  14'd798,  -14'd655,  -14'd1006,  -14'd411,  14'd24,  14'd409,  -14'd32,  -14'd202,  -14'd1160,  14'd171,  14'd773,  14'd1526,  14'd198,  -14'd865,  
14'd1289,  14'd276,  -14'd1252,  14'd1531,  14'd195,  -14'd226,  -14'd705,  14'd300,  -14'd555,  -14'd613,  14'd1574,  -14'd26,  -14'd429,  -14'd686,  14'd557,  14'd447,  
14'd664,  14'd190,  14'd556,  14'd404,  -14'd1519,  14'd1060,  -14'd190,  14'd860,  -14'd495,  -14'd1685,  14'd1256,  14'd500,  14'd1417,  14'd164,  -14'd966,  14'd1141,  
-14'd373,  14'd1172,  -14'd286,  14'd126,  14'd7,  14'd1751,  14'd1465,  14'd1,  14'd1002,  14'd944,  14'd878,  -14'd925,  14'd312,  14'd1100,  -14'd1415,  14'd649,  
-14'd75,  -14'd573,  -14'd950,  -14'd320,  14'd2014,  -14'd922,  -14'd1402,  -14'd451,  -14'd470,  14'd1038,  14'd1324,  -14'd1672,  -14'd60,  -14'd1051,  14'd554,  -14'd731,  
-14'd1028,  14'd1132,  -14'd142,  -14'd208,  14'd423,  -14'd181,  -14'd1777,  -14'd119,  -14'd276,  -14'd224,  -14'd1059,  -14'd637,  -14'd149,  -14'd1256,  -14'd1008,  14'd1004,  
14'd737,  -14'd757,  -14'd176,  -14'd353,  14'd243,  -14'd825,  14'd236,  -14'd4,  14'd871,  -14'd619,  14'd242,  14'd772,  -14'd1833,  -14'd128,  -14'd67,  14'd897,  
14'd1119,  14'd580,  -14'd724,  -14'd1773,  -14'd708,  14'd215,  14'd667,  -14'd688,  -14'd409,  -14'd946,  14'd130,  14'd870,  -14'd910,  14'd532,  14'd210,  -14'd803,  
-14'd1330,  14'd283,  -14'd1027,  14'd874,  -14'd452,  -14'd886,  -14'd222,  14'd164,  -14'd813,  -14'd1041,  14'd543,  -14'd681,  -14'd468,  14'd758,  14'd270,  -14'd1086,  
-14'd317,  14'd529,  -14'd641,  -14'd521,  14'd1536,  14'd1459,  -14'd88,  -14'd481,  14'd1792,  -14'd951,  14'd1949,  14'd750,  14'd639,  -14'd1293,  14'd1312,  14'd962,  
-14'd492,  -14'd1019,  -14'd963,  -14'd1297,  14'd1623,  -14'd1313,  14'd228,  -14'd1090,  -14'd212,  14'd568,  14'd211,  -14'd803,  -14'd454,  -14'd641,  -14'd343,  -14'd817,  
14'd348,  14'd925,  -14'd255,  -14'd619,  -14'd97,  -14'd394,  -14'd894,  -14'd2101,  14'd1827,  14'd1391,  -14'd230,  14'd1125,  -14'd654,  14'd1976,  14'd121,  -14'd421,  
-14'd266,  14'd422,  -14'd33,  -14'd375,  -14'd776,  -14'd568,  -14'd90,  -14'd1125,  14'd176,  -14'd220,  -14'd66,  14'd178,  14'd123,  14'd1908,  -14'd866,  14'd245,  
-14'd1503,  -14'd221,  14'd1363,  14'd762,  14'd16,  -14'd231,  14'd462,  14'd885,  14'd1218,  -14'd837,  -14'd387,  -14'd1508,  -14'd1384,  -14'd147,  -14'd136,  -14'd1441,  

14'd820,  14'd783,  14'd1301,  -14'd1324,  -14'd343,  14'd707,  14'd816,  14'd202,  14'd1319,  14'd74,  -14'd1379,  -14'd573,  14'd303,  -14'd164,  -14'd450,  14'd569,  
-14'd1100,  14'd1889,  14'd1170,  14'd552,  14'd1519,  14'd133,  -14'd633,  -14'd488,  -14'd1532,  -14'd307,  -14'd2199,  14'd657,  14'd820,  -14'd569,  14'd732,  14'd692,  
14'd815,  -14'd638,  -14'd582,  14'd34,  -14'd776,  -14'd1919,  14'd597,  -14'd500,  14'd457,  14'd214,  14'd24,  14'd628,  -14'd1551,  14'd394,  14'd179,  14'd164,  
-14'd1017,  -14'd1311,  14'd1560,  -14'd394,  -14'd456,  -14'd1321,  -14'd307,  14'd328,  -14'd296,  -14'd1152,  -14'd327,  -14'd920,  -14'd1331,  14'd1779,  14'd506,  14'd979,  
-14'd997,  14'd1524,  14'd596,  14'd51,  -14'd757,  14'd398,  14'd385,  14'd111,  14'd1495,  -14'd336,  -14'd199,  -14'd1428,  -14'd1074,  14'd1645,  -14'd540,  14'd1109,  
14'd255,  14'd774,  -14'd653,  -14'd772,  14'd721,  -14'd361,  14'd179,  14'd1637,  -14'd725,  -14'd456,  -14'd1295,  -14'd31,  -14'd1676,  14'd342,  -14'd1001,  14'd3,  
-14'd879,  -14'd601,  14'd197,  14'd207,  14'd1374,  14'd470,  -14'd1121,  14'd536,  -14'd345,  14'd849,  -14'd2261,  14'd599,  -14'd714,  -14'd1897,  14'd542,  -14'd874,  
-14'd495,  -14'd788,  14'd178,  -14'd462,  14'd43,  14'd717,  -14'd330,  -14'd1095,  14'd355,  14'd1034,  14'd45,  -14'd316,  -14'd742,  -14'd740,  -14'd558,  -14'd979,  
-14'd977,  -14'd1745,  14'd1420,  -14'd160,  -14'd548,  -14'd1114,  -14'd24,  14'd244,  -14'd791,  -14'd377,  14'd675,  14'd181,  -14'd1081,  14'd1125,  14'd990,  -14'd917,  
-14'd1033,  14'd216,  -14'd506,  -14'd430,  -14'd108,  14'd518,  -14'd127,  14'd1996,  -14'd67,  14'd450,  -14'd429,  14'd321,  14'd633,  14'd877,  -14'd1233,  -14'd2151,  
14'd41,  -14'd280,  14'd323,  -14'd640,  14'd1588,  -14'd3,  -14'd1120,  14'd7,  14'd970,  14'd38,  -14'd1440,  14'd381,  14'd1075,  -14'd1187,  -14'd959,  14'd40,  
14'd446,  14'd1454,  14'd999,  14'd761,  -14'd1001,  14'd871,  -14'd837,  14'd525,  -14'd812,  14'd1333,  14'd1515,  14'd712,  14'd960,  -14'd1365,  14'd278,  14'd1549,  
-14'd93,  -14'd1062,  -14'd19,  14'd1324,  14'd454,  14'd1519,  -14'd676,  14'd1927,  -14'd936,  -14'd752,  14'd1851,  14'd897,  14'd1227,  -14'd686,  -14'd603,  -14'd119,  
14'd126,  -14'd544,  -14'd444,  -14'd775,  -14'd906,  -14'd1107,  14'd1082,  -14'd1410,  14'd1413,  -14'd300,  14'd1610,  -14'd74,  14'd443,  -14'd19,  -14'd774,  -14'd581,  
14'd664,  -14'd630,  -14'd2163,  14'd1088,  -14'd400,  14'd890,  14'd49,  14'd829,  14'd467,  -14'd717,  -14'd227,  14'd261,  14'd1187,  -14'd1015,  14'd764,  14'd1062,  
14'd197,  -14'd1429,  -14'd1270,  14'd374,  14'd405,  14'd166,  14'd1144,  14'd722,  14'd16,  14'd221,  14'd2545,  14'd204,  14'd1570,  14'd1533,  14'd1205,  14'd521,  
14'd1018,  -14'd1506,  14'd1331,  14'd473,  14'd341,  14'd1114,  14'd548,  -14'd255,  -14'd960,  14'd461,  -14'd163,  -14'd169,  14'd1357,  14'd227,  14'd648,  14'd769,  
14'd31,  14'd1463,  14'd1462,  14'd1088,  14'd300,  14'd510,  -14'd46,  -14'd837,  -14'd413,  -14'd294,  14'd1380,  14'd63,  -14'd980,  -14'd844,  -14'd737,  14'd991,  
14'd127,  14'd732,  14'd291,  14'd242,  14'd1875,  14'd200,  -14'd328,  -14'd61,  -14'd477,  -14'd464,  14'd582,  14'd122,  14'd290,  14'd184,  -14'd747,  -14'd892,  
14'd1387,  -14'd293,  -14'd395,  14'd1525,  -14'd1415,  14'd846,  14'd161,  -14'd153,  14'd500,  14'd962,  -14'd84,  14'd328,  -14'd236,  14'd489,  -14'd133,  -14'd1018,  
14'd879,  14'd1011,  14'd1107,  14'd306,  -14'd1305,  -14'd134,  -14'd54,  -14'd25,  -14'd881,  14'd698,  14'd1322,  -14'd1121,  14'd1393,  14'd950,  14'd435,  -14'd145,  
-14'd345,  14'd406,  -14'd869,  -14'd306,  -14'd166,  -14'd441,  14'd1039,  -14'd292,  -14'd641,  -14'd189,  -14'd600,  -14'd111,  14'd1511,  14'd568,  -14'd94,  -14'd363,  
14'd981,  14'd739,  14'd658,  14'd902,  -14'd7,  14'd728,  -14'd640,  -14'd781,  14'd1033,  -14'd692,  14'd593,  -14'd542,  -14'd340,  -14'd379,  -14'd517,  -14'd149,  
-14'd1395,  14'd1595,  14'd914,  -14'd178,  -14'd860,  -14'd393,  -14'd693,  14'd946,  14'd900,  -14'd61,  -14'd716,  -14'd22,  -14'd295,  14'd960,  14'd951,  14'd1694,  
14'd1780,  14'd202,  14'd1694,  14'd736,  14'd405,  -14'd248,  14'd837,  14'd1060,  14'd1271,  14'd266,  14'd537,  14'd1546,  -14'd650,  14'd184,  14'd1692,  14'd810,  

14'd77,  14'd414,  14'd1900,  -14'd544,  -14'd1862,  -14'd345,  14'd1708,  -14'd854,  -14'd529,  -14'd1614,  14'd463,  -14'd507,  -14'd1146,  14'd1788,  14'd829,  14'd113,  
-14'd716,  -14'd446,  14'd649,  -14'd11,  14'd1031,  -14'd474,  14'd2131,  -14'd2033,  14'd756,  -14'd733,  14'd2897,  -14'd581,  -14'd802,  14'd406,  -14'd1052,  -14'd969,  
14'd360,  14'd157,  14'd109,  -14'd1687,  -14'd43,  -14'd1563,  -14'd129,  -14'd1738,  14'd980,  14'd707,  14'd873,  14'd479,  14'd704,  14'd2429,  -14'd701,  -14'd1138,  
14'd963,  14'd902,  -14'd1375,  -14'd290,  -14'd1196,  -14'd549,  14'd742,  14'd638,  14'd1223,  -14'd566,  14'd438,  -14'd1306,  -14'd311,  -14'd1350,  -14'd170,  -14'd653,  
14'd1943,  14'd819,  -14'd778,  14'd1838,  -14'd443,  14'd240,  -14'd962,  14'd696,  -14'd163,  -14'd309,  -14'd172,  14'd1291,  14'd1757,  14'd1998,  14'd506,  14'd1775,  
-14'd46,  14'd700,  14'd462,  -14'd904,  14'd21,  14'd443,  14'd1629,  -14'd47,  -14'd1480,  -14'd772,  -14'd767,  14'd1218,  -14'd919,  14'd938,  -14'd387,  -14'd995,  
14'd786,  -14'd1465,  -14'd357,  -14'd240,  -14'd170,  -14'd655,  14'd1227,  14'd578,  14'd902,  -14'd1305,  -14'd372,  14'd1177,  14'd113,  14'd217,  14'd75,  -14'd519,  
-14'd129,  -14'd552,  14'd184,  14'd1122,  14'd512,  -14'd150,  -14'd1105,  -14'd1804,  14'd1246,  14'd2382,  14'd1312,  -14'd57,  -14'd932,  14'd579,  -14'd543,  -14'd813,  
-14'd170,  -14'd785,  -14'd3076,  -14'd1354,  -14'd99,  -14'd579,  -14'd1649,  14'd720,  -14'd111,  14'd979,  14'd317,  -14'd1876,  14'd1293,  -14'd1475,  -14'd935,  14'd512,  
-14'd1554,  -14'd79,  -14'd806,  14'd388,  14'd1087,  14'd1248,  -14'd1323,  -14'd310,  -14'd1211,  14'd1995,  14'd798,  14'd217,  14'd1207,  -14'd1012,  -14'd302,  14'd575,  
14'd151,  -14'd230,  14'd923,  14'd1015,  -14'd624,  -14'd204,  14'd541,  -14'd500,  14'd978,  14'd368,  -14'd362,  14'd248,  14'd790,  14'd1024,  14'd1679,  14'd928,  
14'd417,  -14'd854,  14'd1405,  14'd1826,  -14'd546,  14'd446,  -14'd860,  14'd1952,  -14'd206,  14'd355,  14'd92,  -14'd851,  14'd1760,  14'd1574,  14'd1146,  -14'd1101,  
-14'd415,  -14'd1225,  -14'd457,  14'd705,  14'd1621,  14'd150,  14'd503,  -14'd1409,  -14'd71,  14'd183,  14'd1081,  14'd509,  14'd354,  -14'd1439,  14'd54,  -14'd964,  
-14'd664,  -14'd585,  -14'd2599,  -14'd362,  -14'd69,  14'd573,  -14'd754,  -14'd399,  14'd1039,  -14'd1260,  14'd765,  14'd86,  14'd348,  -14'd1396,  -14'd952,  -14'd503,  
-14'd1728,  14'd15,  -14'd565,  14'd2095,  -14'd194,  14'd493,  -14'd1861,  14'd786,  14'd228,  14'd1060,  14'd1779,  -14'd688,  14'd573,  -14'd165,  14'd433,  -14'd571,  
14'd222,  14'd142,  14'd712,  14'd11,  -14'd37,  14'd890,  14'd353,  -14'd638,  -14'd979,  -14'd42,  -14'd132,  14'd270,  14'd770,  14'd314,  -14'd354,  -14'd244,  
14'd35,  -14'd676,  14'd158,  14'd1032,  14'd1020,  -14'd1295,  -14'd2400,  -14'd379,  -14'd1282,  -14'd203,  -14'd578,  14'd382,  14'd333,  14'd347,  14'd394,  14'd602,  
14'd1315,  14'd245,  14'd1867,  -14'd161,  14'd709,  14'd40,  14'd1266,  -14'd558,  -14'd793,  14'd190,  -14'd217,  14'd1672,  14'd1256,  14'd954,  14'd4,  14'd291,  
14'd259,  -14'd78,  14'd72,  -14'd441,  14'd2243,  14'd97,  14'd200,  -14'd345,  14'd664,  -14'd964,  14'd1640,  14'd1047,  -14'd452,  14'd507,  -14'd114,  -14'd440,  
-14'd6,  14'd758,  14'd398,  -14'd184,  14'd705,  14'd194,  14'd47,  14'd968,  14'd277,  -14'd408,  -14'd749,  -14'd922,  -14'd1715,  14'd829,  -14'd126,  -14'd1114,  
14'd1169,  14'd199,  -14'd481,  -14'd602,  -14'd251,  14'd130,  14'd1330,  14'd124,  14'd1105,  14'd288,  -14'd180,  14'd101,  14'd482,  -14'd278,  -14'd800,  14'd554,  
-14'd732,  -14'd626,  14'd78,  -14'd200,  -14'd714,  -14'd420,  -14'd766,  -14'd918,  14'd959,  14'd502,  14'd1421,  -14'd173,  14'd795,  -14'd2346,  14'd788,  14'd717,  
-14'd770,  14'd361,  14'd1045,  14'd193,  -14'd800,  -14'd1610,  14'd540,  -14'd259,  14'd882,  14'd928,  14'd382,  14'd253,  -14'd350,  14'd1355,  14'd51,  14'd340,  
-14'd1057,  14'd234,  14'd1238,  -14'd677,  -14'd1001,  -14'd400,  -14'd269,  14'd940,  14'd558,  -14'd719,  -14'd1408,  -14'd173,  14'd857,  14'd246,  14'd497,  -14'd454,  
-14'd729,  14'd374,  14'd13,  -14'd116,  -14'd1355,  14'd398,  -14'd660,  14'd943,  -14'd651,  -14'd1508,  -14'd738,  -14'd1249,  -14'd51,  14'd1481,  14'd772,  -14'd1324,  

-14'd2,  14'd678,  -14'd481,  14'd250,  -14'd1522,  -14'd548,  14'd1025,  14'd628,  14'd782,  14'd34,  -14'd529,  -14'd101,  -14'd509,  -14'd664,  14'd1724,  14'd294,  
-14'd163,  14'd631,  -14'd94,  14'd613,  -14'd76,  14'd883,  -14'd699,  14'd980,  14'd818,  14'd819,  14'd1785,  -14'd907,  -14'd1363,  -14'd1897,  14'd463,  14'd386,  
14'd701,  14'd611,  -14'd716,  14'd519,  14'd349,  14'd525,  -14'd2184,  -14'd0,  14'd229,  14'd50,  14'd1374,  -14'd129,  14'd1035,  -14'd2636,  14'd321,  -14'd343,  
14'd66,  -14'd566,  14'd713,  -14'd60,  -14'd842,  14'd731,  -14'd1727,  14'd688,  -14'd172,  14'd288,  -14'd650,  -14'd111,  14'd174,  -14'd3790,  -14'd139,  14'd572,  
-14'd1376,  -14'd1577,  14'd318,  -14'd858,  -14'd400,  -14'd845,  -14'd980,  -14'd102,  14'd552,  14'd535,  -14'd325,  14'd744,  -14'd655,  14'd301,  -14'd655,  14'd31,  
-14'd68,  -14'd974,  14'd2096,  14'd1705,  -14'd369,  14'd500,  -14'd776,  14'd703,  -14'd209,  -14'd66,  14'd262,  14'd682,  14'd805,  -14'd701,  14'd37,  14'd442,  
-14'd1538,  -14'd717,  -14'd299,  -14'd133,  14'd602,  14'd1115,  14'd1149,  14'd482,  14'd458,  -14'd195,  -14'd291,  14'd209,  -14'd803,  -14'd847,  -14'd117,  14'd336,  
-14'd2169,  -14'd257,  -14'd1517,  14'd1438,  14'd700,  14'd1008,  -14'd1709,  -14'd482,  -14'd745,  -14'd213,  -14'd494,  -14'd901,  -14'd940,  -14'd1473,  -14'd320,  -14'd927,  
-14'd1163,  14'd937,  14'd2,  -14'd1211,  14'd1016,  14'd84,  -14'd869,  -14'd1209,  -14'd1445,  14'd1521,  -14'd861,  -14'd1329,  -14'd445,  -14'd642,  14'd199,  14'd616,  
-14'd2551,  -14'd218,  14'd272,  -14'd177,  -14'd710,  -14'd714,  14'd536,  14'd135,  14'd410,  14'd761,  14'd338,  -14'd1816,  -14'd543,  14'd156,  -14'd279,  -14'd1226,  
14'd184,  14'd335,  14'd704,  14'd1035,  14'd842,  14'd430,  -14'd139,  14'd930,  -14'd1873,  14'd10,  14'd649,  14'd965,  14'd1056,  14'd903,  14'd422,  14'd354,  
-14'd1474,  14'd655,  -14'd799,  14'd230,  14'd1740,  -14'd211,  -14'd495,  14'd169,  14'd1893,  14'd316,  14'd986,  14'd895,  14'd198,  -14'd1974,  -14'd235,  -14'd394,  
14'd287,  14'd601,  14'd113,  -14'd439,  14'd1710,  14'd116,  14'd38,  14'd366,  14'd23,  14'd477,  14'd376,  14'd833,  -14'd1227,  14'd773,  -14'd704,  14'd1235,  
14'd746,  -14'd1403,  14'd1398,  -14'd234,  -14'd1182,  -14'd266,  -14'd304,  -14'd84,  -14'd869,  -14'd1848,  14'd741,  -14'd98,  14'd240,  14'd848,  14'd1003,  -14'd324,  
14'd1127,  -14'd1190,  14'd1408,  -14'd1044,  -14'd269,  14'd1653,  -14'd308,  14'd308,  14'd1061,  14'd322,  -14'd166,  -14'd243,  14'd127,  14'd918,  -14'd27,  14'd656,  
14'd2047,  14'd51,  14'd204,  -14'd1162,  -14'd1055,  -14'd565,  14'd871,  -14'd875,  14'd1202,  -14'd92,  14'd998,  14'd1515,  -14'd1144,  -14'd1230,  14'd31,  -14'd917,  
-14'd78,  -14'd331,  -14'd1542,  14'd417,  -14'd198,  -14'd371,  -14'd161,  -14'd1080,  14'd1810,  -14'd540,  14'd89,  14'd1492,  14'd894,  14'd660,  -14'd1231,  14'd1197,  
14'd746,  -14'd674,  -14'd344,  14'd28,  -14'd881,  14'd1105,  14'd1086,  -14'd587,  14'd602,  -14'd388,  -14'd1067,  14'd335,  14'd861,  -14'd551,  -14'd757,  14'd488,  
14'd1166,  14'd690,  14'd1535,  14'd786,  14'd1068,  -14'd717,  14'd149,  14'd466,  -14'd91,  -14'd430,  14'd501,  -14'd1573,  14'd794,  14'd2,  14'd796,  14'd54,  
-14'd1167,  14'd1315,  -14'd948,  -14'd285,  -14'd243,  -14'd1264,  -14'd875,  -14'd267,  -14'd511,  14'd1904,  14'd301,  14'd220,  14'd1484,  -14'd167,  14'd455,  -14'd832,  
14'd1437,  14'd1219,  14'd341,  -14'd357,  14'd434,  -14'd47,  14'd2555,  -14'd373,  -14'd475,  -14'd1577,  14'd327,  14'd1218,  -14'd1004,  -14'd497,  -14'd1416,  14'd600,  
14'd112,  14'd407,  -14'd1407,  -14'd535,  -14'd489,  -14'd268,  14'd2830,  -14'd568,  14'd1547,  14'd583,  14'd603,  -14'd396,  -14'd605,  14'd1134,  -14'd1455,  -14'd1250,  
14'd239,  -14'd547,  14'd906,  -14'd294,  14'd33,  -14'd648,  -14'd204,  -14'd324,  14'd562,  14'd109,  -14'd124,  -14'd1440,  14'd912,  14'd1363,  -14'd570,  -14'd1121,  
-14'd121,  14'd1507,  14'd181,  -14'd492,  -14'd391,  14'd1820,  -14'd334,  14'd443,  -14'd123,  14'd815,  14'd318,  -14'd690,  14'd472,  -14'd797,  14'd75,  14'd387,  
-14'd2185,  -14'd1860,  -14'd1753,  14'd1285,  14'd247,  14'd1130,  14'd539,  -14'd560,  -14'd811,  14'd1361,  -14'd954,  -14'd1533,  -14'd686,  -14'd1551,  14'd1088,  -14'd472,  

14'd1174,  14'd374,  14'd105,  14'd193,  -14'd625,  14'd374,  14'd1763,  14'd429,  14'd437,  -14'd416,  14'd877,  14'd608,  14'd90,  14'd738,  -14'd120,  14'd476,  
14'd512,  14'd739,  14'd1277,  14'd646,  14'd695,  14'd421,  14'd244,  -14'd66,  14'd926,  14'd851,  14'd2057,  14'd252,  14'd291,  14'd1077,  -14'd47,  -14'd736,  
-14'd718,  -14'd1628,  14'd692,  -14'd197,  14'd198,  14'd936,  14'd1406,  14'd1490,  -14'd270,  14'd998,  14'd850,  14'd705,  14'd343,  -14'd663,  14'd867,  14'd642,  
-14'd219,  -14'd845,  14'd742,  14'd590,  -14'd1124,  -14'd193,  -14'd227,  -14'd205,  -14'd499,  14'd1222,  -14'd1244,  -14'd75,  14'd1103,  -14'd369,  -14'd740,  14'd11,  
-14'd618,  -14'd540,  -14'd1286,  -14'd1119,  -14'd50,  -14'd782,  -14'd158,  -14'd69,  -14'd635,  14'd164,  14'd32,  -14'd710,  14'd708,  14'd235,  -14'd478,  -14'd531,  
-14'd41,  14'd985,  -14'd422,  14'd745,  14'd442,  14'd1157,  -14'd508,  -14'd128,  14'd540,  14'd883,  -14'd128,  -14'd757,  -14'd1006,  14'd1301,  14'd148,  -14'd1111,  
-14'd376,  14'd91,  14'd1124,  -14'd1017,  -14'd649,  -14'd1254,  -14'd88,  14'd180,  14'd450,  14'd159,  14'd1028,  14'd112,  -14'd138,  14'd1307,  14'd199,  14'd975,  
-14'd146,  -14'd1396,  14'd56,  14'd555,  -14'd240,  14'd843,  -14'd111,  14'd445,  14'd18,  14'd377,  -14'd1195,  -14'd529,  14'd1070,  14'd842,  14'd335,  14'd432,  
-14'd487,  -14'd1799,  14'd6,  14'd702,  14'd804,  14'd547,  -14'd194,  14'd480,  -14'd264,  -14'd737,  -14'd536,  -14'd1195,  -14'd256,  14'd102,  -14'd210,  14'd46,  
-14'd3235,  -14'd1176,  -14'd1617,  -14'd651,  -14'd1097,  -14'd2366,  -14'd118,  -14'd325,  -14'd1990,  -14'd209,  -14'd105,  14'd577,  -14'd1745,  14'd635,  -14'd936,  -14'd529,  
-14'd1430,  -14'd1568,  14'd1487,  -14'd308,  14'd546,  14'd581,  -14'd761,  14'd1173,  14'd685,  14'd1376,  -14'd1467,  -14'd266,  14'd98,  14'd2290,  14'd1021,  -14'd207,  
14'd63,  -14'd443,  14'd706,  14'd976,  -14'd205,  -14'd384,  -14'd1347,  -14'd189,  -14'd1412,  -14'd1661,  -14'd138,  14'd19,  14'd458,  14'd62,  14'd1575,  14'd383,  
14'd93,  -14'd393,  14'd966,  14'd807,  -14'd1214,  14'd517,  -14'd1955,  -14'd726,  14'd752,  14'd602,  -14'd445,  -14'd961,  14'd110,  -14'd952,  14'd204,  -14'd133,  
14'd387,  -14'd833,  -14'd335,  -14'd691,  -14'd235,  14'd666,  -14'd775,  -14'd903,  -14'd1017,  -14'd616,  -14'd1159,  -14'd540,  -14'd988,  14'd472,  14'd197,  -14'd1483,  
-14'd15,  -14'd577,  14'd140,  14'd134,  -14'd1270,  14'd303,  14'd261,  14'd299,  14'd302,  14'd1218,  -14'd563,  14'd206,  -14'd1642,  -14'd585,  -14'd1265,  14'd395,  
-14'd1632,  14'd463,  -14'd588,  -14'd217,  14'd1410,  14'd462,  -14'd1386,  14'd1359,  14'd113,  14'd1387,  -14'd1480,  -14'd133,  14'd149,  14'd242,  -14'd1195,  -14'd864,  
-14'd964,  14'd1356,  14'd652,  -14'd271,  -14'd1183,  14'd104,  -14'd2136,  14'd58,  14'd528,  -14'd484,  14'd1023,  14'd246,  -14'd1103,  -14'd803,  -14'd301,  -14'd376,  
-14'd1319,  -14'd337,  14'd151,  -14'd1294,  14'd65,  -14'd1693,  14'd837,  14'd433,  -14'd1731,  -14'd319,  -14'd583,  14'd938,  14'd474,  14'd126,  -14'd362,  14'd1385,  
14'd348,  14'd356,  14'd79,  14'd242,  -14'd1180,  -14'd576,  14'd74,  14'd45,  14'd1214,  14'd178,  -14'd449,  14'd1651,  14'd114,  14'd1018,  14'd1534,  -14'd345,  
-14'd886,  14'd428,  14'd705,  -14'd1570,  -14'd1369,  14'd582,  14'd1408,  14'd584,  -14'd1120,  14'd1294,  14'd12,  14'd28,  -14'd643,  -14'd722,  14'd865,  -14'd1624,  
-14'd1999,  14'd376,  -14'd1654,  14'd504,  14'd1688,  -14'd1225,  14'd894,  -14'd581,  14'd2143,  -14'd303,  -14'd34,  -14'd662,  -14'd653,  -14'd624,  -14'd366,  -14'd465,  
-14'd45,  -14'd449,  -14'd1361,  -14'd309,  14'd1792,  14'd878,  14'd346,  -14'd1874,  14'd661,  14'd495,  14'd1118,  14'd110,  -14'd624,  -14'd1627,  -14'd39,  14'd1083,  
14'd1025,  14'd1115,  -14'd330,  14'd0,  -14'd549,  -14'd688,  -14'd346,  -14'd635,  14'd1002,  14'd322,  14'd496,  14'd872,  14'd423,  14'd665,  -14'd314,  -14'd949,  
14'd1225,  14'd689,  14'd856,  14'd494,  14'd1182,  14'd2053,  14'd734,  14'd974,  -14'd458,  14'd346,  -14'd172,  14'd990,  14'd1658,  -14'd13,  14'd23,  14'd774,  
14'd851,  -14'd576,  14'd1515,  -14'd24,  14'd332,  14'd631,  14'd1247,  14'd972,  14'd310,  -14'd1198,  -14'd15,  14'd1500,  14'd332,  14'd11,  14'd124,  -14'd347,  

14'd1721,  14'd159,  14'd1813,  14'd538,  14'd28,  14'd895,  14'd351,  -14'd1684,  -14'd355,  14'd543,  14'd611,  14'd607,  -14'd287,  -14'd761,  14'd276,  -14'd149,  
-14'd88,  14'd817,  14'd1557,  -14'd29,  -14'd24,  14'd731,  -14'd276,  -14'd459,  14'd80,  -14'd779,  -14'd780,  14'd394,  -14'd366,  -14'd267,  -14'd11,  14'd595,  
14'd202,  14'd173,  -14'd1299,  14'd546,  14'd310,  14'd126,  14'd278,  14'd866,  14'd1021,  -14'd454,  14'd274,  14'd77,  -14'd1298,  14'd373,  -14'd712,  14'd595,  
14'd165,  -14'd620,  14'd588,  -14'd1896,  14'd270,  -14'd166,  14'd371,  -14'd480,  14'd1354,  14'd138,  14'd276,  14'd1397,  -14'd1310,  14'd3020,  -14'd1045,  -14'd1055,  
-14'd412,  14'd320,  14'd1099,  14'd692,  14'd35,  14'd285,  14'd307,  -14'd59,  14'd833,  -14'd127,  -14'd94,  -14'd277,  -14'd829,  14'd1933,  -14'd947,  -14'd536,  
-14'd247,  14'd1263,  -14'd735,  -14'd602,  -14'd522,  14'd1330,  14'd616,  -14'd277,  -14'd217,  14'd31,  14'd159,  -14'd230,  -14'd616,  14'd259,  14'd320,  14'd111,  
-14'd45,  -14'd322,  14'd1367,  -14'd1261,  -14'd217,  14'd1147,  14'd295,  14'd845,  -14'd580,  14'd42,  -14'd959,  -14'd50,  -14'd539,  14'd894,  14'd1911,  -14'd534,  
14'd2420,  -14'd1168,  14'd1661,  14'd763,  14'd756,  14'd37,  14'd1467,  -14'd242,  -14'd201,  14'd143,  -14'd405,  14'd1128,  -14'd440,  -14'd8,  14'd367,  -14'd1645,  
-14'd157,  -14'd1233,  -14'd139,  14'd949,  14'd614,  14'd75,  14'd552,  -14'd1339,  14'd259,  -14'd418,  -14'd1644,  14'd38,  14'd1221,  14'd1545,  -14'd791,  -14'd414,  
14'd366,  -14'd115,  -14'd723,  14'd711,  14'd1827,  14'd1256,  14'd1076,  14'd350,  14'd762,  -14'd659,  -14'd879,  -14'd964,  14'd204,  14'd1528,  -14'd2038,  -14'd669,  
-14'd331,  14'd1517,  14'd10,  14'd225,  14'd113,  -14'd378,  14'd1373,  14'd329,  -14'd704,  -14'd535,  14'd64,  -14'd1035,  14'd452,  -14'd350,  -14'd761,  14'd1012,  
-14'd421,  -14'd722,  14'd655,  14'd956,  14'd1537,  14'd1469,  14'd1114,  14'd715,  14'd480,  -14'd1101,  -14'd1340,  -14'd1205,  14'd857,  14'd1017,  -14'd933,  14'd48,  
14'd1334,  14'd817,  -14'd433,  -14'd102,  -14'd68,  14'd1695,  -14'd773,  14'd385,  14'd848,  -14'd1333,  -14'd751,  14'd385,  14'd699,  -14'd1609,  14'd1675,  -14'd1340,  
14'd130,  -14'd158,  14'd276,  -14'd489,  -14'd15,  14'd178,  14'd305,  -14'd916,  -14'd631,  14'd322,  -14'd298,  14'd132,  -14'd66,  14'd425,  14'd1036,  14'd695,  
14'd642,  -14'd1903,  -14'd710,  -14'd359,  14'd1467,  14'd588,  14'd1387,  14'd429,  -14'd609,  14'd588,  -14'd1179,  -14'd1019,  -14'd167,  14'd1906,  14'd197,  14'd369,  
14'd1148,  14'd750,  14'd681,  14'd805,  -14'd1306,  -14'd445,  14'd832,  14'd581,  14'd264,  -14'd38,  -14'd56,  -14'd56,  -14'd179,  14'd793,  -14'd577,  14'd641,  
14'd1169,  -14'd281,  14'd195,  14'd522,  14'd2506,  -14'd354,  14'd716,  14'd529,  14'd1259,  14'd47,  -14'd752,  -14'd621,  -14'd43,  14'd1811,  -14'd382,  14'd226,  
14'd221,  14'd418,  -14'd207,  14'd64,  14'd701,  14'd64,  -14'd647,  -14'd917,  -14'd479,  -14'd865,  -14'd1488,  14'd227,  -14'd1322,  14'd1364,  -14'd87,  14'd709,  
-14'd2,  -14'd1598,  14'd823,  -14'd705,  -14'd547,  14'd228,  14'd43,  14'd268,  14'd1061,  -14'd1340,  -14'd918,  14'd628,  -14'd630,  -14'd246,  14'd601,  14'd384,  
-14'd1304,  14'd105,  -14'd66,  14'd99,  -14'd880,  14'd16,  14'd1866,  14'd23,  14'd1224,  -14'd1528,  -14'd156,  -14'd546,  -14'd123,  -14'd1223,  -14'd11,  14'd350,  
14'd510,  14'd127,  -14'd273,  14'd701,  -14'd37,  -14'd1379,  -14'd1487,  -14'd241,  -14'd1259,  14'd594,  -14'd2038,  -14'd1289,  14'd9,  14'd1178,  -14'd121,  14'd367,  
-14'd539,  14'd1541,  14'd263,  14'd563,  14'd725,  -14'd403,  -14'd852,  14'd220,  -14'd1109,  14'd46,  -14'd1556,  -14'd767,  -14'd258,  14'd1343,  14'd1197,  14'd225,  
14'd932,  14'd1078,  14'd370,  -14'd1152,  -14'd181,  14'd200,  14'd71,  14'd922,  -14'd27,  -14'd984,  -14'd1044,  -14'd1041,  -14'd925,  14'd1748,  14'd2388,  -14'd691,  
14'd531,  -14'd848,  14'd459,  14'd93,  14'd1136,  -14'd754,  14'd1194,  14'd1209,  -14'd547,  -14'd1869,  -14'd682,  -14'd995,  14'd591,  14'd2219,  14'd761,  14'd1405,  
14'd172,  14'd1141,  -14'd120,  14'd825,  14'd2116,  14'd1457,  14'd542,  14'd672,  -14'd635,  -14'd1827,  14'd189,  -14'd330,  -14'd759,  14'd1024,  14'd112,  -14'd1062,  

14'd971,  -14'd1008,  -14'd1735,  14'd59,  -14'd405,  14'd64,  -14'd1162,  -14'd68,  -14'd87,  14'd965,  -14'd1786,  -14'd59,  14'd1304,  14'd235,  14'd1680,  14'd557,  
-14'd175,  14'd465,  14'd686,  14'd439,  -14'd376,  14'd49,  -14'd2037,  14'd2077,  14'd890,  14'd1402,  14'd210,  -14'd240,  -14'd338,  -14'd156,  14'd963,  14'd508,  
-14'd15,  -14'd1415,  14'd1004,  14'd310,  -14'd954,  14'd139,  -14'd186,  14'd1056,  14'd436,  14'd116,  14'd3,  14'd1089,  -14'd387,  -14'd480,  14'd1107,  14'd237,  
14'd361,  14'd336,  14'd1653,  14'd385,  -14'd1614,  -14'd1163,  -14'd1765,  14'd72,  14'd151,  14'd876,  -14'd712,  14'd644,  14'd1175,  -14'd1677,  14'd941,  -14'd1075,  
14'd722,  14'd1185,  14'd243,  14'd1027,  -14'd828,  -14'd386,  14'd222,  14'd1200,  14'd192,  14'd788,  -14'd45,  14'd215,  14'd1039,  -14'd1269,  14'd331,  14'd1149,  
14'd97,  14'd1121,  -14'd235,  14'd1615,  14'd218,  14'd972,  -14'd2018,  -14'd1075,  14'd1143,  14'd1682,  -14'd1297,  14'd218,  14'd1000,  -14'd714,  14'd688,  -14'd1097,  
-14'd937,  14'd152,  14'd622,  14'd1370,  -14'd574,  14'd113,  -14'd360,  14'd0,  14'd476,  14'd1599,  -14'd768,  -14'd981,  14'd857,  14'd1646,  14'd663,  14'd294,  
14'd35,  14'd982,  14'd1787,  14'd727,  14'd340,  -14'd1409,  14'd109,  -14'd769,  14'd603,  -14'd113,  14'd1168,  -14'd233,  14'd934,  14'd1927,  -14'd612,  14'd1490,  
-14'd968,  14'd1383,  14'd674,  -14'd437,  -14'd582,  14'd907,  -14'd237,  14'd525,  -14'd1014,  -14'd433,  14'd824,  14'd677,  -14'd213,  14'd359,  14'd281,  -14'd776,  
14'd1354,  -14'd722,  14'd581,  14'd236,  -14'd1263,  14'd955,  14'd480,  14'd645,  -14'd405,  -14'd650,  14'd213,  14'd1703,  14'd404,  -14'd1281,  -14'd567,  -14'd1128,  
-14'd931,  14'd1022,  -14'd67,  14'd125,  14'd1201,  -14'd201,  -14'd1855,  14'd1490,  -14'd1537,  -14'd352,  -14'd391,  14'd229,  -14'd862,  14'd354,  14'd72,  -14'd24,  
14'd99,  14'd631,  14'd309,  -14'd405,  14'd1495,  14'd67,  14'd1435,  -14'd213,  14'd269,  14'd566,  14'd351,  14'd235,  14'd28,  -14'd1119,  -14'd502,  14'd211,  
-14'd957,  -14'd1452,  14'd1332,  -14'd1133,  14'd937,  14'd884,  14'd572,  14'd321,  14'd226,  14'd357,  14'd644,  14'd681,  -14'd1680,  14'd1999,  14'd72,  -14'd1229,  
14'd449,  -14'd764,  -14'd608,  14'd1450,  14'd677,  -14'd1632,  -14'd194,  14'd1339,  14'd355,  14'd81,  -14'd514,  -14'd675,  -14'd0,  -14'd288,  14'd448,  -14'd108,  
14'd1869,  14'd1544,  14'd23,  -14'd927,  14'd56,  -14'd1158,  -14'd203,  14'd579,  -14'd185,  -14'd1630,  -14'd1011,  -14'd387,  -14'd183,  14'd168,  14'd1454,  14'd843,  
14'd681,  -14'd709,  -14'd386,  -14'd574,  -14'd355,  -14'd1909,  14'd606,  -14'd1290,  14'd496,  -14'd451,  -14'd957,  14'd1860,  14'd387,  -14'd831,  -14'd761,  -14'd76,  
14'd1590,  14'd714,  14'd272,  -14'd70,  -14'd297,  14'd272,  14'd3620,  -14'd603,  14'd2481,  -14'd98,  14'd582,  14'd72,  14'd832,  14'd1896,  -14'd127,  14'd541,  
-14'd857,  14'd360,  -14'd232,  14'd255,  14'd303,  14'd1104,  -14'd179,  -14'd776,  14'd952,  -14'd1051,  14'd501,  -14'd609,  -14'd41,  14'd135,  -14'd707,  14'd418,  
-14'd1463,  -14'd182,  -14'd837,  14'd426,  -14'd223,  -14'd1119,  14'd648,  -14'd1851,  14'd320,  14'd1589,  -14'd775,  -14'd1813,  -14'd1024,  -14'd947,  -14'd141,  -14'd1343,  
-14'd788,  14'd51,  -14'd199,  -14'd181,  14'd302,  -14'd576,  14'd170,  -14'd238,  -14'd526,  14'd1427,  -14'd136,  14'd192,  -14'd822,  -14'd1463,  14'd148,  14'd1226,  
14'd396,  -14'd344,  14'd1813,  -14'd490,  -14'd619,  -14'd431,  14'd1462,  14'd57,  14'd337,  14'd571,  -14'd14,  -14'd761,  14'd998,  14'd2024,  -14'd732,  14'd561,  
-14'd174,  14'd206,  14'd676,  14'd637,  -14'd415,  14'd375,  -14'd859,  14'd849,  -14'd1958,  -14'd746,  -14'd542,  -14'd142,  -14'd50,  14'd1686,  -14'd106,  14'd201,  
14'd1246,  -14'd1197,  -14'd908,  -14'd1199,  -14'd1304,  -14'd1121,  -14'd1580,  14'd224,  -14'd1811,  -14'd1350,  14'd821,  -14'd359,  -14'd316,  -14'd50,  14'd347,  14'd1341,  
14'd1619,  14'd508,  -14'd1009,  -14'd161,  -14'd1625,  -14'd481,  -14'd911,  14'd697,  -14'd382,  -14'd468,  14'd151,  -14'd204,  14'd693,  14'd543,  14'd72,  14'd629,  
14'd22,  14'd1058,  14'd2068,  -14'd1421,  14'd245,  -14'd318,  14'd497,  -14'd5,  -14'd299,  -14'd1818,  -14'd328,  -14'd216,  -14'd268,  -14'd423,  -14'd643,  14'd443,  

-14'd487,  -14'd1820,  -14'd472,  14'd878,  14'd1698,  -14'd505,  -14'd1871,  -14'd683,  14'd23,  14'd1132,  -14'd1488,  14'd918,  14'd481,  -14'd1692,  14'd658,  -14'd1091,  
14'd1234,  -14'd1450,  -14'd497,  -14'd337,  14'd1587,  14'd49,  -14'd448,  14'd79,  -14'd769,  14'd151,  -14'd603,  -14'd144,  14'd526,  14'd612,  14'd659,  -14'd776,  
14'd783,  -14'd164,  14'd1574,  14'd425,  -14'd823,  -14'd220,  -14'd189,  14'd14,  14'd330,  -14'd624,  -14'd878,  14'd1691,  -14'd1110,  14'd212,  14'd996,  -14'd707,  
14'd462,  14'd121,  14'd1061,  14'd963,  -14'd344,  14'd287,  14'd459,  14'd1166,  -14'd671,  -14'd882,  -14'd115,  14'd411,  -14'd389,  14'd1,  14'd857,  -14'd559,  
14'd1336,  14'd208,  14'd565,  14'd2186,  -14'd115,  14'd171,  -14'd102,  -14'd793,  14'd1377,  -14'd274,  -14'd438,  14'd532,  -14'd82,  -14'd1937,  14'd1630,  -14'd899,  
-14'd135,  14'd155,  14'd669,  14'd1842,  -14'd1215,  14'd1310,  14'd234,  -14'd530,  -14'd217,  14'd2,  -14'd919,  14'd1281,  -14'd885,  14'd967,  14'd69,  -14'd162,  
14'd893,  -14'd1852,  -14'd1365,  14'd210,  -14'd871,  14'd935,  14'd142,  14'd842,  14'd769,  14'd677,  14'd129,  14'd58,  -14'd320,  -14'd555,  14'd690,  14'd1046,  
-14'd550,  -14'd668,  -14'd292,  14'd1061,  -14'd181,  -14'd657,  14'd52,  14'd119,  -14'd820,  14'd58,  -14'd1143,  -14'd100,  -14'd778,  14'd2204,  14'd174,  -14'd303,  
14'd250,  14'd176,  -14'd194,  -14'd578,  -14'd167,  -14'd215,  -14'd749,  14'd1930,  -14'd2006,  -14'd1332,  -14'd1005,  14'd418,  14'd76,  14'd361,  14'd1931,  -14'd347,  
14'd1811,  14'd2366,  14'd1804,  -14'd706,  -14'd1253,  -14'd96,  14'd278,  -14'd808,  14'd253,  -14'd1992,  -14'd698,  14'd183,  -14'd1793,  -14'd12,  14'd1863,  14'd427,  
-14'd694,  14'd1155,  14'd1168,  14'd273,  14'd295,  -14'd62,  14'd2019,  -14'd248,  14'd1344,  14'd538,  -14'd635,  -14'd935,  -14'd297,  -14'd313,  14'd719,  14'd485,  
14'd108,  -14'd1751,  -14'd626,  -14'd967,  14'd1296,  -14'd746,  14'd1962,  -14'd527,  -14'd42,  -14'd964,  -14'd312,  14'd957,  14'd1190,  14'd1536,  14'd165,  14'd136,  
-14'd1479,  14'd1025,  14'd419,  -14'd642,  -14'd649,  -14'd1345,  -14'd728,  14'd1859,  -14'd2162,  14'd682,  -14'd107,  -14'd665,  -14'd850,  14'd504,  14'd545,  -14'd60,  
-14'd475,  -14'd69,  14'd1707,  -14'd866,  -14'd1280,  14'd87,  -14'd728,  14'd1685,  14'd238,  -14'd1740,  -14'd90,  14'd504,  -14'd1977,  14'd182,  14'd1617,  -14'd209,  
14'd219,  -14'd17,  14'd1821,  14'd242,  -14'd1080,  -14'd882,  -14'd765,  14'd1047,  14'd179,  -14'd1215,  -14'd1407,  14'd636,  -14'd1143,  -14'd614,  14'd377,  -14'd444,  
14'd14,  14'd194,  -14'd652,  -14'd101,  -14'd225,  14'd1131,  14'd1886,  14'd536,  -14'd1255,  -14'd243,  -14'd200,  -14'd829,  14'd218,  -14'd359,  14'd678,  14'd1204,  
14'd564,  -14'd78,  14'd158,  14'd1496,  14'd1180,  -14'd265,  -14'd337,  14'd951,  -14'd659,  -14'd1043,  -14'd845,  -14'd820,  14'd369,  -14'd1402,  14'd353,  -14'd1118,  
-14'd1119,  14'd149,  -14'd228,  -14'd849,  -14'd321,  -14'd1753,  -14'd838,  14'd888,  -14'd1405,  14'd997,  -14'd37,  -14'd1747,  14'd230,  14'd1136,  14'd16,  -14'd1528,  
14'd73,  14'd51,  14'd1533,  14'd167,  14'd747,  14'd932,  14'd1134,  -14'd654,  14'd464,  -14'd1151,  14'd365,  14'd1364,  14'd257,  -14'd687,  -14'd829,  -14'd493,  
14'd2263,  14'd268,  14'd1363,  -14'd116,  -14'd1371,  14'd1256,  14'd548,  14'd859,  -14'd1343,  -14'd443,  -14'd991,  -14'd136,  14'd261,  -14'd1130,  -14'd226,  14'd1122,  
14'd1360,  14'd892,  14'd994,  14'd586,  14'd441,  14'd855,  -14'd703,  14'd1706,  -14'd1033,  14'd530,  14'd157,  -14'd773,  14'd713,  14'd1526,  14'd756,  -14'd83,  
-14'd788,  14'd118,  14'd1788,  14'd390,  14'd99,  14'd432,  -14'd96,  14'd298,  14'd337,  14'd771,  -14'd796,  14'd565,  14'd183,  14'd1197,  -14'd220,  -14'd1077,  
-14'd1392,  -14'd1315,  -14'd129,  14'd163,  -14'd1035,  -14'd369,  14'd1268,  -14'd30,  -14'd1047,  -14'd1338,  -14'd423,  14'd355,  14'd99,  -14'd269,  14'd1057,  14'd218,  
-14'd203,  14'd396,  -14'd34,  -14'd158,  14'd778,  -14'd1491,  14'd506,  -14'd774,  -14'd401,  14'd2007,  14'd676,  -14'd667,  -14'd639,  -14'd605,  -14'd719,  -14'd663,  
14'd760,  14'd437,  -14'd411,  14'd139,  14'd760,  -14'd701,  14'd329,  14'd1587,  -14'd1018,  -14'd1033,  -14'd251,  14'd554,  -14'd745,  14'd901,  -14'd1085,  14'd167,  

-14'd381,  14'd362,  -14'd1079,  -14'd823,  14'd750,  14'd297,  14'd582,  -14'd118,  -14'd328,  14'd335,  14'd649,  14'd613,  -14'd216,  14'd1272,  -14'd712,  -14'd566,  
14'd1102,  -14'd503,  14'd75,  -14'd464,  -14'd924,  14'd53,  -14'd954,  -14'd294,  14'd974,  -14'd1086,  -14'd778,  -14'd159,  -14'd0,  -14'd445,  -14'd1325,  14'd8,  
14'd19,  -14'd305,  -14'd1172,  -14'd294,  -14'd651,  14'd152,  -14'd1515,  14'd140,  -14'd1003,  14'd424,  -14'd959,  -14'd172,  14'd979,  -14'd1775,  -14'd103,  14'd942,  
-14'd156,  14'd81,  -14'd1005,  -14'd729,  -14'd538,  -14'd374,  14'd680,  -14'd475,  -14'd404,  -14'd1607,  14'd310,  -14'd1384,  14'd618,  -14'd1126,  -14'd257,  -14'd795,  
-14'd1779,  14'd358,  -14'd1165,  14'd116,  14'd163,  14'd223,  14'd815,  14'd677,  14'd414,  14'd561,  -14'd356,  14'd378,  -14'd651,  -14'd1391,  14'd917,  -14'd297,  
-14'd1277,  -14'd777,  -14'd808,  -14'd905,  -14'd424,  14'd1396,  14'd975,  -14'd35,  -14'd694,  14'd406,  -14'd54,  14'd73,  -14'd1041,  14'd141,  -14'd1246,  14'd871,  
14'd433,  -14'd1397,  -14'd85,  -14'd438,  -14'd1193,  -14'd628,  -14'd223,  14'd682,  -14'd35,  -14'd1290,  -14'd947,  -14'd387,  -14'd508,  -14'd903,  14'd257,  14'd299,  
14'd496,  14'd1077,  -14'd340,  -14'd503,  14'd1119,  -14'd314,  -14'd144,  -14'd1429,  14'd104,  -14'd123,  14'd226,  14'd159,  -14'd847,  -14'd105,  -14'd352,  -14'd449,  
-14'd459,  -14'd1088,  -14'd1634,  -14'd692,  -14'd1203,  14'd1308,  14'd213,  -14'd830,  14'd211,  14'd636,  -14'd8,  -14'd71,  -14'd1835,  -14'd1215,  -14'd1115,  14'd676,  
14'd327,  -14'd848,  -14'd124,  -14'd1079,  -14'd559,  14'd976,  -14'd155,  14'd200,  14'd670,  14'd1004,  -14'd210,  -14'd55,  14'd545,  -14'd83,  -14'd264,  14'd806,  
-14'd261,  -14'd446,  14'd464,  14'd969,  14'd30,  -14'd861,  -14'd240,  -14'd65,  -14'd1672,  14'd669,  -14'd243,  -14'd654,  -14'd314,  14'd278,  14'd654,  14'd294,  
-14'd809,  -14'd631,  -14'd295,  14'd341,  -14'd386,  14'd695,  14'd43,  -14'd1589,  14'd209,  14'd493,  -14'd552,  14'd1204,  -14'd542,  14'd947,  -14'd205,  14'd247,  
14'd165,  -14'd134,  14'd399,  -14'd253,  14'd9,  -14'd1381,  -14'd392,  -14'd742,  -14'd230,  -14'd305,  -14'd251,  14'd227,  -14'd174,  -14'd1068,  14'd100,  14'd862,  
14'd595,  -14'd828,  14'd220,  14'd591,  14'd835,  14'd112,  -14'd937,  -14'd396,  -14'd107,  -14'd600,  -14'd976,  -14'd130,  -14'd1214,  14'd1222,  14'd730,  -14'd493,  
14'd359,  -14'd98,  -14'd891,  -14'd993,  -14'd978,  -14'd828,  14'd399,  -14'd717,  14'd1031,  -14'd771,  14'd644,  -14'd672,  14'd99,  14'd76,  14'd1044,  14'd541,  
-14'd295,  -14'd413,  -14'd1485,  14'd434,  -14'd174,  -14'd810,  -14'd1737,  14'd447,  -14'd562,  14'd482,  -14'd1469,  -14'd748,  -14'd693,  14'd568,  -14'd1048,  -14'd301,  
-14'd561,  -14'd756,  14'd927,  14'd182,  -14'd452,  14'd231,  -14'd48,  -14'd312,  14'd187,  14'd291,  -14'd1552,  14'd18,  -14'd910,  -14'd1123,  14'd613,  -14'd957,  
-14'd626,  -14'd885,  -14'd1077,  14'd467,  -14'd1258,  14'd119,  -14'd374,  14'd846,  -14'd1109,  -14'd563,  -14'd721,  14'd123,  -14'd1061,  14'd315,  -14'd1346,  14'd637,  
14'd625,  14'd285,  -14'd209,  14'd318,  -14'd20,  -14'd220,  14'd601,  -14'd559,  -14'd893,  -14'd476,  -14'd40,  -14'd447,  14'd680,  -14'd702,  -14'd828,  14'd112,  
14'd259,  14'd455,  -14'd200,  14'd692,  -14'd791,  -14'd11,  -14'd1450,  -14'd115,  -14'd1574,  14'd672,  -14'd902,  -14'd373,  14'd547,  -14'd614,  14'd1492,  14'd1310,  
14'd989,  -14'd701,  14'd287,  -14'd853,  -14'd691,  -14'd221,  14'd659,  -14'd802,  -14'd586,  -14'd720,  14'd1028,  14'd1148,  -14'd620,  -14'd1302,  -14'd1233,  14'd387,  
-14'd342,  14'd1065,  -14'd633,  -14'd443,  -14'd381,  14'd178,  -14'd946,  -14'd41,  -14'd847,  14'd574,  -14'd152,  14'd20,  -14'd339,  -14'd1573,  -14'd964,  -14'd1469,  
14'd1230,  -14'd76,  14'd1108,  -14'd808,  -14'd393,  14'd376,  -14'd460,  -14'd950,  -14'd538,  -14'd51,  -14'd1099,  -14'd584,  -14'd123,  14'd76,  -14'd54,  14'd192,  
-14'd833,  14'd405,  -14'd309,  14'd1423,  -14'd1489,  -14'd878,  -14'd380,  14'd432,  14'd892,  -14'd69,  -14'd621,  -14'd1358,  14'd91,  -14'd1071,  14'd1111,  14'd516,  
14'd799,  14'd1236,  14'd519,  14'd255,  -14'd765,  -14'd356,  -14'd565,  14'd277,  -14'd781,  -14'd6,  -14'd215,  -14'd672,  14'd933,  14'd554,  14'd896,  -14'd390,  

-14'd961,  -14'd1390,  -14'd1254,  -14'd447,  -14'd95,  -14'd463,  -14'd2029,  14'd762,  14'd894,  14'd1698,  14'd670,  -14'd106,  14'd1158,  14'd596,  14'd828,  -14'd77,  
-14'd1126,  14'd945,  14'd156,  14'd961,  -14'd522,  -14'd329,  -14'd1352,  14'd1174,  14'd49,  14'd983,  -14'd370,  -14'd21,  14'd580,  -14'd819,  14'd1372,  -14'd774,  
-14'd669,  14'd640,  14'd1141,  14'd1667,  -14'd911,  14'd826,  -14'd69,  14'd475,  -14'd480,  -14'd1431,  -14'd1174,  14'd820,  14'd1333,  -14'd2101,  14'd1286,  14'd820,  
-14'd418,  -14'd959,  14'd194,  14'd911,  14'd256,  -14'd618,  -14'd1599,  14'd1192,  -14'd660,  14'd1480,  14'd329,  14'd237,  -14'd1101,  -14'd2850,  14'd2194,  -14'd246,  
14'd879,  -14'd487,  14'd434,  14'd381,  -14'd308,  14'd804,  14'd570,  14'd887,  14'd1196,  14'd1292,  14'd520,  14'd139,  -14'd138,  -14'd330,  14'd443,  -14'd820,  
14'd480,  14'd1382,  14'd1161,  14'd312,  -14'd983,  14'd1776,  -14'd57,  -14'd9,  14'd570,  -14'd1023,  -14'd762,  14'd481,  14'd1194,  -14'd87,  14'd145,  -14'd349,  
14'd1228,  -14'd769,  14'd18,  -14'd320,  14'd47,  -14'd99,  -14'd623,  14'd621,  14'd794,  -14'd1632,  -14'd419,  14'd927,  14'd597,  14'd1432,  -14'd248,  14'd865,  
-14'd378,  14'd1179,  14'd12,  -14'd1232,  -14'd730,  14'd1613,  14'd18,  -14'd326,  -14'd73,  -14'd631,  -14'd913,  -14'd602,  -14'd835,  14'd281,  14'd276,  14'd310,  
-14'd613,  14'd1258,  14'd206,  -14'd298,  -14'd670,  14'd145,  -14'd955,  14'd348,  -14'd151,  14'd1013,  -14'd130,  -14'd986,  -14'd509,  14'd1013,  14'd714,  14'd1051,  
-14'd945,  -14'd721,  -14'd713,  14'd366,  14'd537,  -14'd787,  14'd665,  -14'd762,  -14'd775,  14'd104,  -14'd89,  14'd358,  -14'd909,  -14'd1265,  14'd691,  14'd967,  
14'd923,  -14'd253,  -14'd454,  14'd685,  14'd35,  14'd88,  -14'd779,  14'd1079,  14'd1464,  14'd610,  -14'd2311,  -14'd269,  -14'd57,  14'd472,  14'd839,  -14'd104,  
14'd1062,  -14'd435,  -14'd657,  -14'd1333,  14'd513,  14'd856,  14'd979,  14'd208,  14'd663,  -14'd1390,  -14'd813,  14'd176,  14'd1633,  14'd391,  14'd910,  14'd1082,  
-14'd958,  14'd1729,  -14'd998,  -14'd1451,  14'd520,  -14'd389,  14'd1155,  -14'd305,  14'd398,  14'd922,  14'd448,  -14'd792,  14'd334,  14'd1387,  -14'd281,  14'd401,  
14'd293,  14'd444,  14'd1123,  14'd844,  -14'd75,  -14'd456,  -14'd98,  14'd289,  -14'd1130,  -14'd717,  14'd202,  14'd328,  -14'd481,  14'd1350,  14'd685,  14'd538,  
14'd186,  -14'd263,  14'd2331,  -14'd777,  -14'd720,  14'd760,  14'd1045,  -14'd1169,  -14'd900,  -14'd702,  -14'd427,  14'd483,  -14'd1563,  -14'd948,  14'd589,  14'd1015,  
14'd275,  14'd323,  -14'd419,  14'd90,  14'd926,  14'd438,  14'd10,  -14'd687,  -14'd1043,  14'd710,  -14'd2118,  -14'd369,  14'd488,  14'd385,  -14'd183,  -14'd572,  
14'd243,  14'd712,  14'd477,  14'd358,  14'd1373,  -14'd64,  14'd506,  14'd1056,  -14'd52,  14'd388,  14'd1114,  -14'd1006,  14'd755,  -14'd982,  -14'd345,  14'd116,  
-14'd890,  14'd1011,  -14'd399,  -14'd306,  -14'd886,  14'd535,  -14'd425,  -14'd528,  14'd754,  -14'd148,  -14'd941,  -14'd255,  -14'd357,  -14'd434,  -14'd334,  14'd335,  
14'd1843,  14'd799,  14'd840,  14'd336,  14'd378,  14'd1484,  -14'd66,  14'd57,  14'd1071,  -14'd799,  14'd1065,  14'd1680,  14'd530,  -14'd902,  -14'd690,  -14'd276,  
14'd524,  14'd1380,  -14'd318,  14'd55,  -14'd488,  -14'd212,  14'd507,  14'd390,  -14'd489,  -14'd62,  14'd80,  -14'd596,  14'd1864,  -14'd467,  -14'd568,  14'd264,  
-14'd840,  14'd823,  -14'd579,  -14'd545,  -14'd303,  -14'd200,  -14'd1005,  -14'd201,  -14'd95,  -14'd467,  -14'd494,  14'd925,  -14'd896,  -14'd541,  -14'd1134,  -14'd215,  
-14'd37,  14'd136,  -14'd532,  14'd878,  14'd249,  14'd83,  14'd856,  -14'd688,  14'd23,  -14'd455,  14'd392,  14'd1311,  -14'd1004,  -14'd1024,  -14'd449,  14'd1525,  
-14'd1444,  -14'd1672,  14'd56,  -14'd1156,  -14'd393,  -14'd154,  14'd663,  -14'd754,  -14'd1239,  14'd735,  -14'd913,  14'd757,  14'd50,  -14'd622,  14'd217,  -14'd869,  
14'd1360,  -14'd878,  14'd655,  -14'd477,  -14'd164,  -14'd749,  14'd677,  -14'd365,  -14'd487,  14'd755,  14'd265,  -14'd1434,  14'd404,  14'd2123,  -14'd1882,  14'd777,  
-14'd985,  -14'd1201,  -14'd331,  -14'd683,  14'd156,  -14'd540,  14'd687,  -14'd662,  -14'd428,  -14'd2398,  -14'd1897,  -14'd705,  14'd519,  -14'd669,  -14'd1676,  14'd536,  

14'd651,  14'd467,  -14'd912,  14'd831,  14'd695,  14'd356,  14'd456,  -14'd372,  14'd277,  -14'd1398,  14'd3018,  14'd338,  -14'd565,  -14'd747,  -14'd749,  -14'd1867,  
-14'd1473,  -14'd1100,  -14'd1341,  14'd730,  -14'd1261,  -14'd921,  -14'd2092,  -14'd1363,  14'd714,  -14'd582,  14'd1117,  14'd433,  -14'd1092,  -14'd805,  -14'd1106,  -14'd915,  
14'd399,  14'd446,  -14'd438,  14'd874,  -14'd88,  14'd1620,  -14'd1771,  14'd1477,  14'd295,  14'd250,  14'd125,  -14'd61,  -14'd886,  -14'd2837,  -14'd860,  14'd1369,  
-14'd1731,  -14'd1249,  14'd1010,  -14'd1326,  -14'd1000,  14'd10,  -14'd88,  -14'd608,  14'd1713,  14'd1418,  14'd250,  -14'd682,  14'd807,  -14'd2052,  -14'd130,  14'd288,  
-14'd433,  -14'd1878,  14'd1687,  -14'd218,  -14'd198,  -14'd1414,  -14'd68,  14'd266,  14'd366,  14'd875,  14'd378,  -14'd812,  -14'd1252,  -14'd362,  -14'd2045,  14'd195,  
14'd1059,  14'd44,  14'd547,  14'd1339,  14'd321,  14'd1034,  -14'd1434,  14'd260,  14'd1406,  14'd1026,  14'd468,  14'd444,  14'd455,  -14'd161,  14'd98,  14'd136,  
14'd201,  14'd925,  14'd328,  -14'd416,  -14'd998,  14'd37,  -14'd681,  -14'd525,  14'd223,  -14'd130,  -14'd543,  -14'd425,  14'd177,  14'd45,  14'd424,  14'd1215,  
14'd113,  -14'd697,  -14'd120,  14'd1593,  -14'd760,  14'd364,  -14'd1596,  14'd44,  -14'd325,  14'd644,  -14'd473,  14'd328,  -14'd880,  -14'd1123,  14'd953,  14'd176,  
-14'd1425,  14'd304,  -14'd815,  -14'd137,  -14'd684,  -14'd320,  14'd1340,  -14'd691,  14'd1008,  14'd1105,  -14'd1009,  -14'd1407,  14'd333,  14'd174,  -14'd248,  -14'd452,  
-14'd1300,  -14'd329,  -14'd934,  14'd1074,  -14'd155,  -14'd252,  -14'd748,  14'd1052,  -14'd108,  14'd1164,  -14'd211,  -14'd369,  14'd129,  -14'd743,  -14'd1718,  -14'd600,  
14'd355,  -14'd281,  -14'd30,  14'd510,  14'd1332,  14'd481,  14'd217,  14'd1130,  -14'd15,  14'd106,  14'd107,  -14'd634,  14'd610,  14'd393,  14'd873,  -14'd171,  
-14'd1182,  14'd350,  -14'd21,  14'd1449,  14'd1161,  -14'd1414,  -14'd319,  -14'd979,  14'd1570,  -14'd697,  14'd1762,  14'd11,  14'd555,  -14'd667,  14'd334,  14'd385,  
14'd561,  14'd907,  -14'd491,  14'd417,  -14'd205,  -14'd825,  -14'd30,  14'd1057,  -14'd1047,  -14'd122,  14'd1251,  14'd461,  -14'd208,  -14'd1026,  -14'd9,  14'd466,  
14'd1686,  -14'd107,  14'd199,  -14'd1011,  14'd294,  -14'd44,  14'd1183,  14'd683,  -14'd666,  -14'd1818,  14'd1131,  -14'd296,  14'd287,  -14'd991,  14'd711,  14'd346,  
-14'd435,  14'd843,  14'd640,  -14'd274,  14'd1190,  14'd1325,  14'd612,  -14'd293,  -14'd271,  14'd752,  14'd480,  -14'd192,  14'd1202,  14'd77,  -14'd791,  -14'd643,  
-14'd992,  14'd1414,  14'd907,  14'd1082,  14'd2016,  -14'd642,  -14'd1563,  14'd357,  -14'd48,  14'd238,  -14'd559,  -14'd537,  14'd612,  14'd19,  -14'd242,  14'd99,  
-14'd820,  14'd772,  -14'd416,  14'd911,  14'd1195,  -14'd442,  -14'd2019,  14'd539,  14'd1270,  -14'd1486,  14'd277,  -14'd459,  14'd643,  -14'd2052,  14'd577,  -14'd22,  
14'd1211,  -14'd1208,  14'd1155,  -14'd1000,  -14'd1049,  -14'd1226,  -14'd673,  14'd34,  -14'd86,  -14'd75,  -14'd1150,  14'd1492,  -14'd570,  14'd1819,  -14'd1119,  -14'd503,  
14'd1672,  14'd127,  14'd1268,  -14'd838,  -14'd1344,  -14'd439,  14'd1363,  -14'd1070,  14'd791,  -14'd345,  14'd381,  14'd1427,  14'd832,  14'd298,  14'd328,  14'd512,  
-14'd369,  -14'd456,  -14'd1902,  -14'd337,  -14'd376,  -14'd420,  -14'd769,  14'd1293,  -14'd855,  14'd219,  14'd858,  14'd69,  -14'd392,  14'd129,  14'd1192,  14'd1069,  
-14'd1375,  14'd1929,  -14'd870,  -14'd1420,  14'd301,  -14'd1442,  14'd2019,  -14'd1078,  14'd1047,  -14'd103,  -14'd1039,  14'd243,  14'd502,  -14'd987,  -14'd251,  -14'd314,  
-14'd77,  -14'd350,  -14'd975,  -14'd678,  -14'd378,  14'd428,  14'd2135,  14'd580,  14'd737,  -14'd1506,  14'd526,  14'd403,  -14'd69,  -14'd922,  -14'd781,  -14'd1167,  
-14'd1366,  -14'd163,  -14'd248,  14'd168,  -14'd1165,  -14'd968,  14'd983,  -14'd1639,  14'd1566,  14'd666,  14'd1029,  -14'd101,  -14'd424,  14'd1317,  14'd1080,  14'd929,  
-14'd1170,  -14'd763,  -14'd408,  14'd1381,  14'd1423,  -14'd955,  14'd980,  -14'd945,  -14'd177,  14'd337,  -14'd909,  14'd254,  -14'd229,  -14'd740,  14'd222,  -14'd297,  
-14'd1010,  -14'd711,  14'd1066,  -14'd134,  -14'd1136,  14'd883,  14'd107,  -14'd366,  -14'd203,  14'd1752,  -14'd1124,  14'd1071,  -14'd139,  14'd317,  14'd744,  14'd520,  

14'd652,  -14'd615,  14'd1200,  -14'd1000,  -14'd1535,  -14'd772,  14'd395,  14'd3,  -14'd264,  14'd834,  14'd1442,  -14'd676,  -14'd571,  -14'd131,  -14'd38,  -14'd698,  
-14'd1226,  -14'd890,  -14'd2128,  -14'd556,  -14'd346,  14'd292,  14'd593,  14'd707,  14'd1063,  -14'd1175,  14'd614,  14'd1543,  14'd1183,  -14'd1316,  -14'd212,  -14'd166,  
14'd86,  14'd167,  -14'd1526,  14'd800,  14'd1736,  14'd1027,  14'd89,  14'd482,  -14'd1119,  14'd579,  14'd1736,  14'd794,  14'd534,  -14'd836,  -14'd942,  -14'd581,  
14'd1757,  14'd1437,  14'd575,  14'd1420,  -14'd121,  14'd706,  -14'd192,  14'd70,  14'd643,  14'd879,  14'd406,  -14'd92,  -14'd454,  -14'd2196,  14'd53,  14'd865,  
-14'd64,  14'd572,  14'd26,  -14'd486,  14'd812,  14'd926,  14'd798,  14'd1609,  -14'd615,  -14'd362,  14'd183,  -14'd695,  14'd2025,  -14'd654,  -14'd1317,  -14'd1011,  
-14'd787,  -14'd1517,  14'd635,  -14'd944,  14'd289,  -14'd144,  -14'd1352,  -14'd383,  14'd1555,  14'd666,  14'd832,  14'd949,  14'd90,  -14'd959,  14'd966,  -14'd1490,  
14'd1015,  14'd780,  14'd559,  -14'd1470,  -14'd74,  -14'd1509,  14'd612,  -14'd1584,  -14'd1244,  -14'd622,  14'd192,  -14'd260,  14'd521,  -14'd745,  -14'd794,  14'd282,  
-14'd860,  14'd131,  14'd587,  14'd853,  14'd1028,  14'd840,  14'd1652,  -14'd807,  -14'd1306,  14'd199,  14'd969,  14'd919,  -14'd156,  -14'd1473,  14'd1410,  -14'd928,  
14'd842,  14'd380,  -14'd1902,  14'd416,  14'd1801,  14'd231,  14'd264,  14'd64,  14'd161,  -14'd721,  14'd951,  -14'd939,  14'd798,  -14'd902,  14'd1064,  14'd440,  
-14'd3202,  -14'd219,  -14'd2021,  14'd725,  -14'd511,  -14'd1057,  14'd49,  -14'd856,  14'd1071,  14'd1587,  14'd952,  14'd260,  14'd1267,  14'd686,  -14'd46,  14'd1778,  
14'd719,  -14'd166,  14'd484,  14'd1051,  -14'd397,  -14'd114,  14'd1287,  -14'd1056,  -14'd987,  -14'd479,  -14'd1499,  -14'd311,  -14'd368,  14'd361,  14'd1291,  14'd965,  
14'd1347,  -14'd541,  14'd495,  14'd1174,  -14'd1554,  14'd330,  14'd590,  -14'd329,  -14'd322,  -14'd1616,  14'd1800,  14'd322,  14'd576,  -14'd1059,  14'd148,  -14'd1153,  
14'd297,  -14'd1430,  -14'd377,  14'd120,  -14'd542,  -14'd59,  14'd1423,  14'd696,  14'd1157,  14'd422,  14'd1885,  -14'd974,  14'd1273,  -14'd995,  14'd73,  -14'd200,  
14'd213,  14'd47,  -14'd507,  14'd424,  -14'd1322,  14'd112,  -14'd1029,  -14'd476,  14'd1003,  -14'd1113,  14'd520,  14'd253,  14'd183,  -14'd46,  14'd1108,  14'd168,  
-14'd2192,  -14'd985,  -14'd182,  14'd1455,  -14'd412,  14'd301,  -14'd173,  -14'd238,  14'd406,  14'd3069,  14'd1542,  14'd1202,  -14'd1361,  14'd1418,  -14'd145,  -14'd1989,  
14'd56,  14'd565,  -14'd2,  14'd1467,  -14'd219,  14'd520,  -14'd477,  -14'd275,  14'd741,  14'd1041,  14'd927,  14'd1297,  -14'd77,  -14'd955,  -14'd1219,  14'd1664,  
14'd1675,  -14'd1248,  14'd643,  14'd1561,  -14'd461,  14'd683,  14'd2535,  14'd1484,  -14'd261,  -14'd1633,  14'd515,  14'd107,  14'd1392,  -14'd505,  14'd64,  14'd887,  
-14'd950,  14'd1133,  -14'd286,  -14'd757,  -14'd469,  14'd412,  14'd571,  -14'd74,  14'd287,  -14'd180,  -14'd1007,  14'd763,  -14'd561,  -14'd496,  -14'd431,  -14'd448,  
14'd1176,  14'd169,  14'd1382,  -14'd900,  -14'd2043,  -14'd468,  14'd470,  14'd1669,  14'd1396,  14'd265,  14'd266,  -14'd578,  -14'd476,  -14'd411,  14'd158,  14'd857,  
14'd1213,  -14'd354,  -14'd1969,  14'd939,  14'd154,  -14'd1372,  14'd328,  14'd1019,  14'd1593,  14'd416,  14'd455,  14'd593,  -14'd1045,  14'd1143,  14'd398,  -14'd314,  
14'd1206,  14'd691,  -14'd72,  -14'd2468,  -14'd1014,  14'd465,  14'd722,  -14'd68,  -14'd2103,  -14'd329,  14'd822,  14'd732,  -14'd1041,  14'd70,  -14'd1372,  14'd453,  
14'd635,  -14'd426,  14'd2591,  -14'd272,  -14'd115,  -14'd272,  14'd1690,  -14'd1304,  14'd550,  14'd282,  -14'd829,  -14'd1362,  14'd260,  14'd263,  -14'd876,  14'd1342,  
-14'd402,  14'd683,  14'd249,  -14'd1530,  14'd1767,  -14'd509,  14'd1028,  14'd166,  14'd2390,  -14'd171,  -14'd1278,  -14'd2100,  -14'd1205,  14'd2324,  14'd1065,  -14'd1266,  
-14'd218,  -14'd2007,  14'd447,  14'd325,  -14'd453,  -14'd1250,  -14'd1132,  -14'd1785,  14'd1977,  -14'd9,  -14'd1434,  -14'd1573,  -14'd2191,  -14'd316,  -14'd169,  -14'd1141,  
-14'd488,  -14'd1763,  14'd27,  14'd57,  -14'd99,  14'd2229,  14'd32,  -14'd368,  14'd788,  14'd1956,  -14'd946,  -14'd610,  -14'd594,  14'd401,  14'd929,  -14'd134,  

14'd232,  -14'd1483,  -14'd147,  -14'd182,  -14'd224,  14'd351,  -14'd541,  14'd1349,  14'd1775,  -14'd327,  -14'd336,  14'd497,  14'd613,  14'd397,  -14'd1174,  -14'd240,  
14'd387,  14'd620,  14'd444,  -14'd1347,  14'd693,  -14'd28,  14'd95,  14'd1162,  14'd1295,  -14'd106,  14'd1105,  -14'd142,  -14'd35,  -14'd1407,  14'd591,  -14'd864,  
14'd16,  -14'd584,  -14'd248,  14'd501,  14'd268,  14'd656,  -14'd800,  14'd23,  -14'd941,  14'd253,  -14'd404,  -14'd15,  -14'd158,  -14'd354,  14'd99,  -14'd407,  
-14'd129,  -14'd365,  -14'd319,  -14'd372,  -14'd147,  -14'd1155,  14'd619,  14'd615,  14'd293,  -14'd45,  -14'd114,  -14'd24,  -14'd1241,  -14'd157,  -14'd627,  -14'd274,  
-14'd359,  -14'd1249,  14'd1431,  -14'd607,  -14'd458,  -14'd45,  -14'd1459,  -14'd121,  14'd936,  14'd274,  -14'd376,  14'd523,  -14'd118,  -14'd1345,  14'd487,  -14'd77,  
-14'd668,  14'd946,  14'd429,  14'd214,  14'd32,  14'd797,  -14'd868,  -14'd78,  14'd939,  -14'd545,  -14'd581,  -14'd60,  14'd655,  -14'd1457,  14'd1112,  14'd142,  
-14'd345,  14'd222,  14'd1,  -14'd17,  -14'd405,  14'd861,  14'd745,  14'd483,  -14'd325,  -14'd953,  -14'd310,  -14'd777,  -14'd854,  14'd11,  -14'd1170,  14'd1132,  
14'd101,  -14'd756,  14'd1238,  14'd864,  14'd429,  -14'd105,  -14'd1405,  -14'd279,  -14'd1366,  -14'd246,  -14'd317,  -14'd1023,  14'd292,  -14'd898,  14'd664,  -14'd544,  
-14'd827,  -14'd857,  -14'd1444,  14'd321,  -14'd162,  14'd19,  -14'd1149,  14'd421,  -14'd135,  -14'd1321,  14'd60,  -14'd195,  -14'd803,  -14'd292,  -14'd1144,  -14'd1061,  
-14'd106,  -14'd649,  14'd805,  14'd220,  14'd385,  -14'd337,  14'd1,  -14'd12,  -14'd1407,  -14'd1345,  14'd992,  -14'd406,  -14'd322,  14'd1395,  14'd190,  -14'd633,  
-14'd38,  14'd81,  -14'd1298,  -14'd323,  14'd615,  14'd490,  14'd465,  14'd388,  -14'd568,  14'd1315,  14'd550,  -14'd941,  14'd382,  -14'd717,  -14'd211,  -14'd501,  
-14'd903,  14'd1329,  -14'd876,  14'd802,  -14'd931,  14'd12,  -14'd497,  14'd267,  14'd257,  -14'd900,  -14'd751,  14'd701,  -14'd668,  14'd499,  -14'd1749,  -14'd445,  
-14'd738,  -14'd115,  14'd143,  14'd805,  -14'd280,  14'd1532,  -14'd1206,  -14'd710,  -14'd866,  -14'd663,  -14'd17,  14'd542,  14'd192,  -14'd574,  14'd836,  -14'd966,  
14'd21,  14'd415,  -14'd976,  -14'd420,  14'd647,  -14'd660,  -14'd17,  -14'd1193,  -14'd1339,  -14'd1191,  -14'd934,  -14'd1308,  -14'd352,  14'd117,  14'd262,  -14'd658,  
14'd890,  14'd241,  14'd1053,  14'd1435,  -14'd1175,  -14'd74,  14'd744,  -14'd581,  -14'd245,  14'd269,  -14'd439,  -14'd565,  14'd529,  -14'd244,  14'd326,  -14'd1455,  
14'd948,  14'd368,  14'd338,  -14'd845,  14'd424,  14'd919,  14'd30,  14'd4,  14'd601,  14'd694,  -14'd418,  -14'd425,  -14'd783,  -14'd940,  -14'd1402,  14'd6,  
14'd15,  -14'd888,  14'd444,  14'd175,  14'd594,  -14'd1616,  -14'd1096,  14'd486,  14'd314,  -14'd13,  14'd597,  -14'd165,  -14'd318,  -14'd957,  -14'd331,  -14'd834,  
14'd50,  -14'd541,  14'd5,  -14'd612,  14'd157,  -14'd415,  -14'd898,  -14'd1284,  -14'd782,  14'd683,  14'd581,  -14'd461,  14'd394,  14'd1317,  14'd235,  -14'd921,  
14'd18,  14'd932,  -14'd609,  -14'd1179,  -14'd1426,  -14'd1170,  -14'd831,  -14'd642,  14'd320,  -14'd399,  14'd64,  -14'd1028,  -14'd532,  14'd400,  -14'd499,  14'd295,  
-14'd1165,  -14'd317,  -14'd132,  -14'd1057,  14'd896,  14'd542,  14'd293,  -14'd503,  -14'd1037,  -14'd793,  -14'd991,  -14'd1154,  -14'd1214,  14'd814,  -14'd162,  -14'd368,  
-14'd1160,  -14'd84,  -14'd979,  14'd206,  14'd87,  14'd354,  -14'd379,  14'd443,  14'd1125,  -14'd214,  14'd1041,  -14'd122,  14'd538,  -14'd1591,  14'd417,  14'd1174,  
-14'd892,  -14'd718,  14'd1346,  14'd392,  14'd34,  14'd1191,  -14'd1227,  -14'd394,  -14'd287,  14'd965,  -14'd812,  14'd590,  -14'd72,  -14'd342,  14'd169,  -14'd361,  
14'd295,  -14'd870,  -14'd487,  -14'd1571,  14'd540,  -14'd809,  14'd591,  14'd16,  -14'd591,  14'd228,  -14'd436,  -14'd329,  14'd161,  -14'd646,  14'd190,  14'd68,  
-14'd704,  -14'd742,  14'd478,  14'd710,  -14'd1080,  -14'd762,  -14'd263,  -14'd1170,  -14'd531,  14'd186,  -14'd1316,  -14'd1313,  14'd118,  -14'd262,  -14'd240,  -14'd91,  
-14'd317,  14'd1352,  14'd1123,  -14'd194,  -14'd1380,  14'd74,  -14'd207,  -14'd689,  -14'd570,  -14'd4,  -14'd1651,  14'd891,  -14'd834,  -14'd817,  -14'd1292,  -14'd53,  

-14'd784,  14'd103,  14'd1669,  14'd1603,  14'd50,  -14'd223,  -14'd1022,  14'd1435,  -14'd205,  14'd864,  14'd120,  -14'd2208,  14'd1147,  14'd820,  -14'd218,  14'd156,  
-14'd1311,  -14'd44,  14'd1816,  14'd787,  -14'd285,  -14'd915,  14'd80,  14'd583,  14'd725,  -14'd10,  14'd257,  -14'd538,  14'd628,  14'd3728,  14'd872,  -14'd329,  
-14'd688,  -14'd370,  14'd2233,  14'd112,  -14'd2036,  -14'd84,  14'd927,  -14'd64,  -14'd257,  14'd771,  -14'd579,  14'd707,  -14'd453,  14'd2886,  14'd246,  -14'd941,  
14'd2059,  14'd551,  14'd889,  -14'd49,  14'd187,  14'd1043,  14'd586,  -14'd1151,  14'd1581,  -14'd53,  14'd1043,  14'd1549,  -14'd918,  -14'd444,  -14'd69,  -14'd1916,  
14'd1892,  14'd2494,  -14'd1817,  14'd1115,  -14'd1299,  14'd832,  14'd1317,  14'd787,  14'd499,  -14'd843,  14'd1372,  -14'd249,  14'd1362,  -14'd1666,  -14'd589,  14'd2026,  
-14'd207,  14'd1113,  -14'd430,  -14'd1320,  14'd2161,  -14'd1138,  -14'd1025,  -14'd655,  -14'd1245,  -14'd1149,  14'd878,  14'd556,  14'd777,  14'd1221,  14'd807,  -14'd806,  
-14'd775,  -14'd224,  14'd1690,  14'd570,  -14'd347,  14'd987,  14'd784,  -14'd1461,  -14'd603,  -14'd172,  14'd113,  14'd314,  14'd133,  14'd1994,  14'd28,  -14'd117,  
-14'd341,  -14'd679,  14'd1682,  14'd1000,  -14'd825,  14'd853,  -14'd39,  -14'd754,  14'd1304,  -14'd1082,  -14'd103,  -14'd982,  -14'd813,  14'd2336,  -14'd559,  -14'd1282,  
14'd283,  -14'd690,  -14'd307,  14'd856,  -14'd793,  -14'd73,  14'd350,  14'd281,  -14'd161,  -14'd929,  -14'd648,  14'd368,  14'd1006,  14'd491,  -14'd718,  -14'd679,  
14'd1398,  -14'd803,  -14'd2359,  14'd645,  14'd331,  -14'd922,  -14'd416,  -14'd614,  14'd1524,  14'd1174,  14'd620,  -14'd850,  -14'd705,  -14'd1501,  -14'd1009,  14'd1034,  
-14'd62,  -14'd1078,  14'd126,  14'd674,  -14'd264,  -14'd1266,  -14'd704,  14'd254,  -14'd948,  -14'd434,  14'd496,  14'd371,  -14'd503,  -14'd624,  14'd756,  -14'd255,  
-14'd514,  -14'd431,  -14'd588,  -14'd751,  -14'd53,  -14'd358,  -14'd92,  -14'd131,  -14'd1085,  -14'd476,  -14'd774,  -14'd643,  -14'd1095,  14'd1811,  -14'd329,  14'd1175,  
14'd385,  -14'd876,  14'd1488,  -14'd1188,  -14'd1258,  14'd880,  -14'd156,  14'd326,  -14'd841,  14'd854,  -14'd1554,  -14'd255,  -14'd487,  14'd905,  14'd142,  14'd257,  
14'd1151,  14'd487,  14'd1561,  14'd1702,  -14'd1265,  14'd1387,  -14'd340,  -14'd637,  14'd796,  -14'd1872,  14'd5,  14'd198,  -14'd1017,  14'd940,  -14'd1281,  -14'd13,  
-14'd622,  -14'd1358,  14'd903,  14'd1213,  -14'd711,  14'd257,  -14'd707,  -14'd529,  14'd883,  -14'd335,  -14'd568,  -14'd1066,  -14'd1930,  -14'd1002,  14'd712,  14'd405,  
-14'd1144,  14'd985,  -14'd1211,  14'd1137,  14'd1189,  14'd399,  14'd1530,  14'd1441,  14'd1327,  14'd339,  14'd908,  -14'd1054,  14'd1038,  -14'd1410,  -14'd1343,  -14'd187,  
-14'd854,  -14'd1270,  14'd547,  14'd228,  -14'd1883,  -14'd1512,  14'd606,  14'd459,  14'd186,  14'd2011,  14'd812,  -14'd482,  14'd316,  -14'd696,  -14'd563,  14'd59,  
14'd333,  -14'd200,  -14'd536,  14'd959,  -14'd83,  14'd344,  14'd217,  14'd24,  -14'd33,  14'd547,  14'd57,  14'd102,  14'd915,  14'd1745,  14'd297,  -14'd1365,  
-14'd1593,  -14'd190,  14'd336,  14'd1300,  -14'd678,  -14'd987,  14'd639,  14'd1348,  -14'd253,  -14'd976,  14'd1350,  -14'd558,  14'd399,  -14'd649,  -14'd1102,  14'd1328,  
14'd736,  -14'd307,  14'd761,  14'd142,  14'd1723,  -14'd447,  14'd346,  14'd87,  -14'd464,  -14'd605,  -14'd447,  14'd1034,  14'd908,  14'd448,  14'd251,  14'd38,  
14'd38,  14'd938,  14'd392,  -14'd1369,  -14'd1504,  -14'd34,  14'd161,  -14'd1161,  -14'd630,  14'd401,  14'd56,  14'd388,  -14'd780,  -14'd855,  14'd181,  14'd1503,  
14'd484,  14'd1009,  14'd1879,  -14'd1723,  14'd413,  14'd129,  14'd1581,  -14'd433,  -14'd69,  14'd288,  14'd391,  14'd452,  14'd1022,  14'd1385,  14'd708,  -14'd77,  
-14'd97,  14'd566,  14'd552,  14'd497,  -14'd1301,  -14'd255,  14'd643,  -14'd1395,  -14'd44,  14'd62,  -14'd1600,  -14'd820,  14'd1338,  14'd1688,  -14'd249,  14'd81,  
-14'd2033,  14'd1084,  -14'd2225,  -14'd383,  14'd462,  -14'd175,  14'd513,  -14'd806,  -14'd847,  -14'd102,  14'd1245,  -14'd2554,  14'd170,  -14'd1119,  14'd733,  14'd681,  
-14'd1584,  14'd171,  -14'd1417,  14'd44,  14'd136,  -14'd191,  -14'd250,  14'd910,  -14'd1643,  -14'd1999,  14'd430,  -14'd2051,  -14'd1221,  14'd1097,  -14'd381,  -14'd276,  

-14'd1937,  -14'd1034,  14'd229,  -14'd791,  14'd2458,  14'd392,  -14'd1219,  14'd1772,  -14'd568,  -14'd281,  14'd533,  -14'd710,  14'd41,  -14'd1950,  -14'd193,  14'd54,  
14'd88,  14'd1586,  14'd837,  -14'd176,  14'd1228,  14'd797,  -14'd168,  14'd1324,  -14'd534,  14'd1317,  -14'd1368,  -14'd938,  14'd1169,  -14'd656,  14'd422,  14'd1120,  
-14'd1093,  -14'd856,  14'd973,  14'd465,  -14'd1102,  14'd672,  14'd99,  -14'd931,  -14'd1797,  14'd189,  -14'd872,  -14'd290,  14'd487,  14'd520,  14'd954,  14'd645,  
-14'd683,  14'd1377,  14'd1225,  14'd343,  14'd115,  14'd667,  14'd323,  14'd316,  14'd1162,  14'd455,  14'd1117,  14'd613,  -14'd1592,  14'd2251,  -14'd1779,  14'd56,  
14'd1859,  14'd1585,  -14'd726,  14'd693,  -14'd7,  14'd988,  14'd1018,  -14'd1183,  14'd1617,  -14'd470,  14'd814,  14'd250,  -14'd496,  14'd934,  14'd689,  14'd1496,  
-14'd1609,  -14'd118,  -14'd2394,  -14'd697,  -14'd664,  -14'd283,  14'd293,  14'd533,  -14'd676,  -14'd126,  14'd1580,  -14'd1293,  -14'd1199,  -14'd1668,  -14'd1006,  14'd472,  
-14'd1466,  -14'd863,  -14'd938,  -14'd658,  14'd1990,  -14'd414,  -14'd1165,  14'd344,  -14'd533,  14'd100,  14'd396,  -14'd653,  -14'd1120,  -14'd1113,  -14'd1021,  -14'd96,  
14'd1150,  -14'd822,  14'd1349,  14'd413,  14'd875,  -14'd493,  14'd471,  -14'd38,  -14'd2183,  14'd846,  -14'd258,  14'd1273,  -14'd118,  -14'd131,  -14'd640,  14'd179,  
14'd1448,  -14'd224,  14'd1808,  14'd559,  14'd1376,  -14'd225,  14'd1055,  14'd571,  14'd507,  -14'd1262,  14'd737,  -14'd408,  14'd459,  14'd1215,  14'd616,  -14'd437,  
14'd1440,  -14'd95,  -14'd17,  14'd760,  -14'd62,  -14'd30,  14'd1370,  14'd289,  14'd723,  14'd545,  -14'd422,  -14'd1196,  14'd568,  -14'd604,  -14'd640,  14'd517,  
-14'd1524,  -14'd1010,  -14'd1871,  -14'd1096,  14'd796,  -14'd1159,  -14'd1155,  14'd555,  14'd1676,  -14'd890,  14'd2238,  -14'd61,  -14'd1143,  -14'd1253,  14'd428,  -14'd1180,  
14'd540,  14'd389,  -14'd345,  14'd525,  -14'd164,  14'd992,  -14'd986,  14'd1008,  -14'd415,  14'd5,  14'd17,  -14'd276,  -14'd839,  14'd710,  14'd764,  14'd238,  
14'd1845,  -14'd850,  -14'd72,  -14'd1327,  14'd268,  -14'd21,  -14'd1046,  14'd866,  14'd707,  14'd1069,  -14'd321,  -14'd277,  14'd1652,  -14'd1561,  -14'd851,  14'd375,  
14'd49,  -14'd1422,  -14'd281,  14'd1196,  14'd970,  -14'd366,  -14'd235,  14'd1239,  -14'd838,  14'd1338,  14'd580,  -14'd467,  14'd1506,  -14'd65,  -14'd1161,  14'd650,  
-14'd1794,  14'd305,  -14'd756,  14'd710,  14'd583,  -14'd1242,  14'd959,  -14'd979,  -14'd1001,  14'd666,  14'd457,  14'd394,  -14'd8,  -14'd1086,  14'd764,  14'd677,  
14'd670,  14'd451,  -14'd1164,  14'd855,  -14'd1092,  -14'd225,  -14'd314,  -14'd735,  14'd948,  -14'd815,  14'd375,  -14'd220,  -14'd782,  14'd1313,  -14'd69,  -14'd876,  
14'd211,  -14'd793,  -14'd94,  14'd905,  -14'd1114,  14'd506,  14'd195,  14'd232,  14'd679,  14'd784,  -14'd547,  -14'd959,  14'd804,  14'd1493,  14'd1532,  -14'd1136,  
-14'd570,  14'd166,  14'd168,  14'd677,  14'd990,  14'd143,  14'd267,  -14'd720,  -14'd370,  -14'd1043,  14'd1278,  14'd1252,  -14'd324,  14'd252,  -14'd800,  14'd1034,  
-14'd259,  -14'd49,  -14'd574,  14'd567,  14'd186,  14'd680,  14'd874,  14'd311,  14'd1045,  14'd1202,  14'd637,  -14'd43,  -14'd1263,  -14'd841,  14'd1196,  14'd748,  
14'd456,  -14'd1899,  -14'd1363,  14'd256,  14'd1033,  -14'd530,  -14'd808,  14'd441,  -14'd673,  14'd753,  14'd2209,  14'd1007,  14'd453,  14'd37,  -14'd597,  14'd1516,  
14'd670,  -14'd138,  14'd1461,  14'd1445,  -14'd378,  -14'd173,  -14'd300,  -14'd418,  14'd873,  14'd80,  -14'd213,  -14'd54,  14'd367,  -14'd317,  14'd446,  14'd897,  
-14'd1064,  -14'd568,  -14'd159,  14'd1751,  14'd111,  14'd1175,  -14'd1049,  -14'd672,  -14'd1192,  14'd1013,  -14'd326,  -14'd244,  14'd325,  14'd1192,  14'd1221,  14'd433,  
14'd594,  14'd561,  14'd346,  -14'd86,  14'd279,  -14'd813,  -14'd1030,  -14'd482,  -14'd1008,  -14'd875,  -14'd211,  -14'd353,  14'd1396,  -14'd535,  14'd621,  14'd1297,  
-14'd104,  14'd1133,  14'd448,  -14'd286,  -14'd708,  14'd55,  -14'd615,  -14'd845,  -14'd891,  -14'd1209,  14'd1182,  14'd98,  14'd737,  14'd494,  -14'd304,  14'd148,  
-14'd151,  14'd2046,  14'd497,  -14'd912,  14'd1035,  14'd84,  -14'd745,  14'd972,  -14'd822,  -14'd447,  14'd31,  -14'd228,  -14'd451,  14'd884,  -14'd207,  14'd362,  

-14'd549,  -14'd1028,  -14'd1175,  -14'd707,  14'd1264,  14'd318,  14'd474,  14'd1045,  -14'd979,  14'd840,  14'd1102,  -14'd165,  14'd2763,  -14'd399,  -14'd161,  -14'd1177,  
14'd990,  -14'd380,  14'd34,  14'd866,  14'd166,  14'd870,  -14'd214,  14'd1027,  -14'd912,  -14'd124,  14'd1016,  14'd816,  14'd57,  14'd260,  14'd820,  14'd994,  
14'd1951,  14'd535,  14'd500,  14'd742,  -14'd279,  14'd183,  -14'd608,  14'd490,  -14'd944,  -14'd1435,  14'd708,  14'd47,  14'd554,  14'd404,  -14'd107,  14'd3,  
14'd136,  14'd507,  -14'd715,  14'd905,  -14'd241,  -14'd72,  -14'd5,  -14'd917,  -14'd1028,  -14'd759,  14'd2233,  -14'd69,  14'd1466,  -14'd296,  -14'd358,  14'd103,  
-14'd179,  -14'd1200,  -14'd1385,  14'd1566,  14'd926,  14'd463,  -14'd432,  14'd1023,  -14'd248,  -14'd1111,  14'd884,  -14'd977,  14'd1010,  14'd1188,  -14'd76,  -14'd664,  
14'd772,  14'd791,  -14'd1062,  -14'd90,  14'd1290,  -14'd529,  -14'd52,  -14'd252,  -14'd892,  -14'd747,  14'd1380,  -14'd1066,  14'd1126,  -14'd866,  14'd46,  -14'd586,  
-14'd722,  14'd371,  -14'd745,  14'd471,  -14'd113,  14'd206,  14'd251,  14'd950,  -14'd825,  -14'd548,  14'd1060,  -14'd1599,  -14'd504,  -14'd1078,  14'd36,  -14'd98,  
-14'd373,  14'd368,  14'd1028,  14'd340,  14'd1111,  14'd632,  -14'd289,  14'd689,  -14'd838,  14'd36,  14'd1514,  -14'd799,  14'd889,  14'd2602,  -14'd557,  14'd1482,  
-14'd1318,  14'd493,  14'd28,  -14'd49,  14'd110,  -14'd290,  -14'd152,  14'd1131,  14'd1270,  14'd582,  14'd1605,  -14'd911,  -14'd194,  14'd241,  14'd821,  14'd549,  
14'd315,  14'd136,  14'd1185,  -14'd229,  14'd390,  -14'd608,  14'd1555,  14'd9,  14'd537,  -14'd283,  14'd1834,  14'd1443,  14'd178,  14'd495,  14'd225,  14'd349,  
-14'd1284,  14'd1809,  -14'd710,  -14'd966,  14'd606,  -14'd1809,  -14'd384,  14'd283,  14'd1647,  14'd309,  14'd2382,  -14'd1012,  14'd122,  14'd3,  -14'd265,  -14'd832,  
-14'd1005,  -14'd540,  -14'd142,  -14'd930,  14'd820,  14'd270,  -14'd1293,  -14'd60,  14'd301,  14'd1672,  -14'd846,  -14'd367,  -14'd1829,  -14'd1255,  -14'd1014,  -14'd170,  
14'd227,  -14'd210,  14'd408,  -14'd1414,  14'd1301,  14'd353,  -14'd384,  14'd70,  14'd723,  14'd1720,  14'd493,  14'd1389,  14'd745,  -14'd66,  14'd572,  14'd471,  
14'd754,  14'd261,  14'd536,  14'd393,  14'd892,  14'd646,  14'd239,  -14'd290,  14'd1633,  -14'd391,  14'd283,  14'd1426,  -14'd406,  14'd790,  14'd1457,  14'd169,  
-14'd1653,  14'd136,  -14'd1701,  14'd265,  -14'd322,  -14'd2322,  14'd83,  -14'd369,  14'd353,  14'd443,  -14'd58,  -14'd792,  14'd878,  14'd373,  14'd1179,  -14'd624,  
14'd269,  -14'd1346,  -14'd179,  -14'd99,  -14'd2016,  14'd332,  -14'd221,  -14'd299,  14'd639,  -14'd1258,  -14'd448,  -14'd376,  14'd298,  -14'd372,  -14'd923,  -14'd160,  
-14'd864,  -14'd1390,  -14'd1050,  14'd653,  -14'd1747,  14'd435,  14'd638,  14'd770,  14'd980,  14'd1170,  14'd434,  14'd1632,  -14'd535,  14'd1042,  14'd823,  -14'd1296,  
-14'd416,  -14'd99,  14'd554,  14'd312,  14'd720,  14'd853,  14'd435,  -14'd48,  -14'd109,  -14'd576,  14'd1078,  14'd284,  14'd914,  -14'd999,  14'd1993,  -14'd1520,  
-14'd1132,  -14'd734,  14'd137,  14'd201,  14'd357,  14'd652,  14'd156,  -14'd39,  14'd430,  14'd153,  -14'd483,  -14'd163,  14'd295,  -14'd860,  -14'd80,  -14'd932,  
14'd133,  14'd612,  -14'd11,  -14'd420,  14'd508,  14'd185,  -14'd720,  14'd402,  -14'd348,  14'd920,  14'd105,  -14'd346,  -14'd1323,  -14'd1042,  -14'd1013,  14'd790,  
-14'd337,  14'd345,  14'd248,  14'd372,  -14'd2075,  14'd451,  -14'd38,  14'd107,  14'd2136,  14'd447,  14'd428,  14'd395,  -14'd1038,  14'd521,  14'd1048,  -14'd298,  
14'd270,  -14'd1091,  14'd20,  14'd862,  14'd565,  -14'd859,  -14'd148,  14'd842,  14'd818,  14'd625,  14'd1148,  14'd579,  -14'd149,  14'd361,  -14'd116,  -14'd281,  
14'd1248,  -14'd1392,  -14'd1016,  14'd610,  -14'd68,  14'd1307,  14'd1261,  14'd1225,  14'd480,  14'd570,  -14'd719,  14'd173,  14'd911,  -14'd1640,  14'd964,  14'd1370,  
14'd101,  14'd1456,  14'd415,  -14'd1068,  14'd856,  -14'd372,  14'd226,  14'd50,  -14'd13,  14'd708,  14'd62,  -14'd389,  -14'd749,  14'd658,  -14'd582,  -14'd318,  
14'd1079,  -14'd1053,  14'd1137,  14'd199,  -14'd1567,  14'd950,  -14'd235,  14'd518,  14'd1042,  14'd2438,  -14'd552,  14'd586,  -14'd471,  14'd41,  -14'd887,  14'd1163,  

14'd950,  -14'd1415,  -14'd793,  -14'd489,  -14'd1499,  14'd501,  14'd1921,  -14'd1418,  14'd997,  -14'd437,  -14'd197,  14'd1141,  -14'd517,  -14'd91,  -14'd1559,  -14'd1616,  
-14'd940,  -14'd833,  -14'd1899,  -14'd117,  -14'd2,  14'd645,  -14'd246,  -14'd683,  -14'd525,  14'd948,  -14'd875,  -14'd375,  -14'd1159,  -14'd253,  14'd403,  -14'd137,  
-14'd1113,  14'd242,  -14'd1343,  -14'd610,  14'd1816,  -14'd572,  -14'd1771,  -14'd237,  -14'd128,  14'd283,  -14'd17,  -14'd679,  -14'd89,  -14'd3548,  -14'd225,  14'd817,  
-14'd1022,  -14'd830,  -14'd1165,  -14'd64,  14'd567,  -14'd135,  -14'd1482,  14'd652,  14'd649,  14'd823,  -14'd1454,  14'd415,  -14'd777,  -14'd396,  -14'd863,  14'd371,  
-14'd1484,  -14'd1229,  14'd989,  14'd99,  -14'd66,  -14'd156,  -14'd789,  -14'd563,  -14'd280,  14'd922,  -14'd1095,  -14'd584,  14'd1411,  -14'd31,  14'd653,  14'd327,  
14'd37,  14'd483,  -14'd388,  -14'd480,  -14'd2219,  14'd279,  14'd209,  14'd857,  14'd375,  14'd409,  14'd1396,  -14'd93,  -14'd8,  -14'd463,  -14'd246,  14'd912,  
14'd728,  14'd691,  -14'd711,  -14'd659,  -14'd1017,  14'd212,  14'd624,  -14'd400,  -14'd191,  14'd522,  -14'd1064,  14'd578,  -14'd958,  14'd956,  14'd413,  14'd1315,  
14'd919,  -14'd1024,  -14'd1642,  -14'd139,  14'd282,  14'd664,  14'd196,  -14'd174,  -14'd140,  14'd102,  -14'd756,  14'd141,  14'd1281,  -14'd2077,  14'd1033,  -14'd154,  
-14'd21,  -14'd930,  -14'd1653,  -14'd90,  14'd300,  -14'd888,  14'd684,  -14'd258,  14'd420,  -14'd860,  14'd464,  14'd111,  14'd625,  -14'd205,  -14'd293,  14'd649,  
-14'd1745,  14'd244,  14'd1517,  14'd81,  14'd89,  -14'd324,  14'd14,  14'd286,  -14'd1102,  -14'd521,  14'd1010,  -14'd1060,  14'd440,  -14'd322,  14'd449,  -14'd469,  
-14'd491,  -14'd62,  14'd804,  14'd369,  14'd487,  -14'd258,  -14'd1846,  14'd1973,  14'd961,  -14'd290,  -14'd3609,  -14'd895,  14'd904,  14'd1406,  14'd1215,  -14'd401,  
14'd226,  14'd660,  -14'd746,  14'd1589,  14'd912,  14'd158,  -14'd1088,  14'd665,  -14'd1347,  -14'd690,  14'd839,  -14'd1045,  14'd1049,  14'd83,  14'd1132,  -14'd590,  
14'd468,  14'd1327,  -14'd1739,  -14'd1268,  14'd104,  14'd830,  14'd1202,  -14'd592,  -14'd516,  -14'd658,  -14'd639,  14'd791,  -14'd127,  -14'd2274,  -14'd884,  -14'd107,  
-14'd811,  14'd665,  14'd490,  -14'd2376,  14'd930,  14'd399,  -14'd705,  14'd136,  -14'd317,  -14'd1218,  -14'd182,  14'd306,  14'd32,  -14'd244,  -14'd1018,  14'd1290,  
14'd680,  14'd7,  14'd96,  -14'd1001,  -14'd889,  14'd1249,  -14'd425,  -14'd550,  14'd1106,  14'd947,  14'd981,  -14'd274,  -14'd1443,  14'd508,  -14'd19,  14'd702,  
-14'd128,  -14'd1760,  -14'd540,  14'd1747,  14'd1309,  14'd1028,  -14'd2169,  14'd182,  -14'd468,  -14'd93,  -14'd684,  14'd67,  14'd974,  14'd247,  14'd6,  -14'd503,  
-14'd305,  -14'd616,  -14'd105,  -14'd121,  14'd2277,  14'd306,  -14'd241,  -14'd489,  14'd121,  -14'd1248,  14'd931,  -14'd262,  14'd1149,  -14'd114,  -14'd171,  14'd13,  
14'd1133,  14'd1893,  14'd316,  -14'd192,  14'd1826,  -14'd1130,  14'd79,  14'd142,  -14'd1345,  -14'd105,  14'd1597,  -14'd954,  -14'd1007,  14'd322,  -14'd948,  -14'd518,  
14'd641,  14'd1104,  -14'd1483,  -14'd555,  14'd1577,  14'd1243,  -14'd431,  -14'd427,  14'd1273,  -14'd384,  -14'd1019,  14'd1317,  -14'd305,  14'd320,  -14'd944,  -14'd1441,  
-14'd1319,  -14'd2061,  14'd398,  -14'd827,  -14'd1301,  14'd218,  -14'd233,  14'd263,  14'd1448,  -14'd12,  -14'd580,  -14'd1477,  14'd1029,  14'd697,  -14'd344,  -14'd1409,  
14'd11,  14'd939,  -14'd336,  14'd1271,  14'd1704,  14'd769,  -14'd197,  14'd32,  14'd528,  14'd1317,  14'd172,  14'd988,  14'd398,  -14'd1476,  14'd1796,  14'd178,  
14'd151,  -14'd506,  14'd396,  14'd1054,  14'd982,  -14'd1483,  14'd356,  -14'd166,  14'd1029,  -14'd1395,  14'd678,  14'd120,  14'd274,  -14'd896,  14'd49,  -14'd703,  
14'd1239,  14'd74,  14'd801,  14'd1028,  14'd171,  14'd1226,  -14'd238,  -14'd508,  14'd1739,  14'd630,  14'd949,  14'd1200,  -14'd14,  -14'd1227,  -14'd683,  14'd323,  
14'd1004,  14'd648,  -14'd90,  -14'd429,  14'd314,  -14'd414,  -14'd454,  -14'd638,  14'd1389,  -14'd504,  -14'd862,  14'd768,  14'd1199,  14'd194,  14'd770,  -14'd664,  
14'd2065,  -14'd1038,  14'd1482,  14'd547,  -14'd969,  14'd798,  14'd1793,  -14'd586,  14'd2871,  14'd644,  -14'd261,  14'd2110,  14'd212,  14'd694,  14'd329,  -14'd845,  

-14'd885,  14'd836,  14'd1113,  -14'd613,  14'd449,  14'd164,  14'd460,  14'd1477,  14'd652,  -14'd526,  -14'd562,  14'd71,  14'd158,  14'd947,  -14'd1082,  14'd1934,  
-14'd275,  14'd1053,  14'd1902,  -14'd2251,  14'd273,  -14'd925,  14'd1483,  14'd462,  -14'd763,  -14'd64,  14'd8,  14'd611,  14'd300,  14'd1034,  14'd130,  -14'd606,  
-14'd845,  14'd103,  14'd496,  -14'd740,  14'd949,  -14'd1589,  14'd792,  -14'd892,  -14'd140,  -14'd584,  14'd1190,  14'd1601,  14'd1364,  14'd3083,  -14'd891,  14'd826,  
-14'd483,  14'd1524,  14'd405,  -14'd642,  14'd1278,  -14'd19,  14'd1720,  14'd765,  -14'd115,  -14'd2191,  -14'd485,  -14'd91,  14'd483,  14'd3436,  -14'd623,  -14'd244,  
14'd949,  14'd410,  -14'd777,  -14'd282,  -14'd1851,  14'd99,  14'd693,  -14'd569,  -14'd540,  -14'd655,  14'd231,  14'd505,  14'd1137,  -14'd22,  -14'd568,  -14'd1005,  
-14'd827,  -14'd260,  -14'd453,  14'd194,  14'd1042,  -14'd840,  14'd104,  -14'd756,  -14'd1066,  14'd878,  -14'd211,  -14'd968,  14'd140,  14'd1536,  14'd575,  -14'd433,  
14'd1209,  -14'd1352,  14'd568,  14'd1734,  -14'd597,  -14'd2,  14'd885,  -14'd48,  -14'd141,  -14'd761,  14'd1071,  14'd506,  -14'd683,  14'd579,  -14'd950,  -14'd914,  
14'd1463,  -14'd1191,  14'd34,  14'd1776,  -14'd73,  -14'd634,  14'd2075,  -14'd777,  -14'd1431,  -14'd120,  -14'd267,  14'd345,  -14'd573,  -14'd1311,  -14'd1359,  -14'd2375,  
14'd2022,  14'd1418,  14'd1303,  -14'd659,  -14'd33,  14'd276,  -14'd152,  -14'd119,  14'd1331,  14'd913,  -14'd510,  14'd352,  14'd435,  14'd585,  -14'd503,  -14'd1164,  
14'd2310,  -14'd595,  -14'd640,  -14'd431,  14'd459,  -14'd155,  14'd1008,  -14'd91,  14'd461,  14'd1151,  -14'd158,  14'd1052,  -14'd591,  -14'd189,  14'd146,  14'd364,  
-14'd700,  14'd196,  14'd902,  -14'd497,  14'd286,  14'd151,  14'd728,  14'd463,  -14'd78,  14'd256,  14'd610,  -14'd1056,  -14'd600,  -14'd1151,  -14'd873,  14'd1540,  
14'd793,  14'd962,  -14'd260,  14'd1422,  -14'd286,  -14'd630,  -14'd609,  14'd145,  -14'd671,  14'd650,  14'd624,  14'd417,  -14'd62,  14'd590,  14'd297,  -14'd241,  
-14'd145,  -14'd1515,  -14'd703,  14'd219,  -14'd180,  14'd881,  -14'd760,  -14'd295,  -14'd221,  14'd220,  14'd280,  -14'd211,  -14'd99,  -14'd1580,  -14'd351,  14'd1009,  
-14'd381,  -14'd225,  14'd135,  14'd994,  14'd405,  14'd320,  -14'd23,  -14'd1282,  14'd675,  14'd117,  -14'd1,  14'd1272,  14'd117,  -14'd527,  -14'd73,  14'd1591,  
-14'd724,  -14'd1144,  14'd325,  14'd123,  14'd222,  14'd725,  -14'd573,  -14'd652,  14'd535,  14'd461,  14'd541,  14'd821,  -14'd325,  -14'd1713,  14'd1941,  14'd624,  
14'd458,  14'd1204,  -14'd495,  -14'd477,  -14'd1568,  -14'd362,  -14'd184,  -14'd123,  -14'd524,  -14'd335,  14'd792,  -14'd431,  14'd1268,  -14'd103,  -14'd82,  14'd598,  
14'd121,  -14'd593,  14'd273,  14'd583,  14'd378,  14'd420,  -14'd395,  -14'd169,  -14'd251,  -14'd692,  -14'd1692,  14'd1000,  -14'd88,  -14'd472,  14'd475,  14'd169,  
14'd97,  14'd862,  -14'd492,  -14'd203,  14'd1399,  14'd184,  -14'd691,  14'd1066,  14'd250,  -14'd589,  14'd450,  14'd427,  -14'd834,  -14'd146,  -14'd742,  -14'd937,  
-14'd29,  -14'd383,  -14'd375,  14'd838,  -14'd427,  14'd570,  14'd1194,  14'd194,  14'd242,  14'd5,  14'd654,  -14'd84,  14'd778,  -14'd664,  -14'd400,  14'd368,  
-14'd610,  14'd2316,  -14'd101,  14'd555,  14'd917,  -14'd340,  14'd376,  -14'd31,  -14'd829,  -14'd1143,  14'd393,  -14'd200,  -14'd85,  14'd1301,  -14'd1139,  14'd116,  
-14'd226,  14'd488,  14'd655,  -14'd2269,  -14'd2369,  14'd274,  14'd1033,  -14'd664,  14'd630,  14'd370,  -14'd968,  -14'd1027,  14'd202,  14'd1627,  -14'd1059,  -14'd569,  
-14'd500,  14'd669,  14'd790,  -14'd699,  -14'd74,  14'd962,  14'd873,  14'd112,  14'd40,  14'd789,  -14'd884,  14'd1642,  -14'd470,  14'd1295,  -14'd412,  14'd242,  
-14'd608,  14'd872,  14'd83,  -14'd749,  -14'd354,  14'd989,  14'd342,  14'd589,  14'd238,  -14'd1286,  -14'd74,  -14'd159,  14'd700,  14'd163,  -14'd84,  -14'd1715,  
-14'd442,  -14'd128,  -14'd1258,  -14'd255,  14'd230,  -14'd458,  14'd843,  -14'd1037,  14'd81,  -14'd190,  14'd62,  -14'd787,  -14'd133,  14'd865,  -14'd179,  14'd737,  
14'd1625,  -14'd1108,  -14'd1226,  -14'd1510,  -14'd1354,  -14'd273,  14'd339,  -14'd354,  -14'd1133,  -14'd2385,  -14'd820,  -14'd2679,  -14'd264,  -14'd380,  -14'd787,  -14'd1650,  

-14'd145,  -14'd759,  14'd295,  14'd250,  -14'd434,  -14'd579,  14'd2341,  -14'd758,  -14'd8,  -14'd91,  -14'd1737,  14'd314,  -14'd2227,  -14'd994,  14'd212,  -14'd29,  
-14'd1687,  -14'd663,  14'd247,  -14'd1105,  -14'd460,  -14'd447,  -14'd327,  -14'd1914,  -14'd1682,  -14'd296,  14'd1014,  -14'd1315,  -14'd644,  14'd59,  -14'd68,  -14'd616,  
-14'd524,  -14'd577,  14'd254,  -14'd1244,  14'd302,  -14'd893,  14'd397,  14'd582,  14'd536,  14'd301,  14'd870,  -14'd511,  14'd358,  -14'd1412,  14'd467,  14'd204,  
-14'd399,  14'd619,  14'd498,  14'd1814,  -14'd507,  14'd1141,  -14'd223,  14'd1167,  14'd983,  -14'd120,  -14'd279,  14'd201,  -14'd362,  14'd259,  -14'd232,  -14'd869,  
14'd434,  14'd334,  -14'd314,  14'd2164,  -14'd1474,  14'd268,  -14'd789,  14'd320,  -14'd462,  -14'd43,  14'd210,  -14'd159,  14'd1883,  14'd4,  14'd737,  -14'd203,  
-14'd255,  -14'd670,  -14'd511,  14'd700,  -14'd1337,  -14'd664,  14'd1134,  -14'd502,  14'd83,  14'd234,  14'd659,  -14'd1207,  14'd160,  -14'd631,  14'd234,  -14'd95,  
14'd1624,  -14'd1156,  -14'd589,  14'd503,  -14'd652,  -14'd1311,  -14'd100,  14'd491,  14'd976,  14'd189,  -14'd527,  -14'd71,  -14'd1216,  14'd697,  14'd142,  -14'd1349,  
-14'd68,  -14'd1932,  -14'd488,  14'd312,  14'd1170,  14'd171,  14'd173,  14'd314,  14'd1817,  14'd1206,  14'd1057,  -14'd693,  14'd355,  -14'd17,  14'd1530,  -14'd609,  
-14'd1198,  14'd366,  -14'd533,  -14'd735,  14'd865,  -14'd1094,  14'd150,  14'd1787,  14'd728,  14'd33,  14'd643,  -14'd1418,  14'd80,  -14'd2032,  14'd153,  14'd867,  
-14'd1897,  -14'd1845,  14'd585,  -14'd394,  14'd772,  14'd90,  -14'd2032,  14'd375,  14'd728,  14'd753,  -14'd0,  14'd70,  14'd1584,  14'd379,  -14'd1448,  -14'd60,  
-14'd286,  14'd457,  -14'd785,  14'd1257,  14'd48,  14'd1043,  -14'd94,  14'd1147,  14'd330,  -14'd409,  -14'd2542,  -14'd867,  14'd66,  14'd1446,  14'd780,  14'd217,  
14'd25,  14'd263,  14'd563,  -14'd79,  -14'd1351,  -14'd579,  -14'd960,  14'd910,  -14'd615,  14'd271,  -14'd325,  -14'd1072,  -14'd663,  14'd671,  14'd400,  -14'd1099,  
-14'd1436,  -14'd96,  -14'd1302,  -14'd23,  14'd704,  14'd616,  -14'd319,  -14'd314,  -14'd864,  14'd206,  14'd388,  -14'd1611,  14'd534,  14'd37,  -14'd1173,  14'd1203,  
-14'd2022,  -14'd719,  -14'd226,  -14'd634,  14'd882,  14'd1040,  -14'd928,  14'd56,  14'd558,  14'd87,  14'd355,  -14'd962,  -14'd44,  -14'd1372,  -14'd598,  14'd1376,  
-14'd2475,  -14'd562,  14'd1526,  14'd873,  14'd758,  -14'd1493,  14'd1021,  -14'd1117,  -14'd761,  14'd896,  -14'd918,  14'd605,  -14'd1613,  14'd210,  14'd757,  -14'd269,  
-14'd450,  14'd715,  14'd265,  14'd1710,  14'd383,  14'd1412,  -14'd441,  -14'd13,  -14'd117,  14'd643,  -14'd115,  -14'd1478,  14'd756,  14'd1466,  -14'd313,  14'd905,  
-14'd795,  14'd873,  -14'd151,  14'd471,  14'd3,  14'd823,  -14'd784,  -14'd497,  -14'd888,  -14'd807,  14'd1176,  -14'd108,  -14'd238,  14'd241,  14'd192,  -14'd157,  
14'd800,  14'd23,  -14'd790,  14'd268,  -14'd805,  -14'd1150,  14'd727,  14'd998,  -14'd1154,  14'd727,  14'd1182,  14'd533,  14'd488,  14'd48,  -14'd459,  -14'd554,  
14'd325,  14'd1798,  -14'd12,  -14'd1743,  14'd151,  14'd635,  14'd581,  14'd700,  14'd1239,  -14'd2308,  -14'd40,  14'd893,  -14'd12,  14'd554,  -14'd614,  14'd476,  
14'd209,  14'd195,  14'd1034,  -14'd958,  14'd627,  -14'd582,  14'd2080,  14'd2277,  -14'd77,  -14'd2255,  -14'd809,  14'd79,  14'd319,  14'd588,  14'd500,  -14'd1326,  
14'd672,  14'd741,  -14'd1609,  14'd592,  14'd2000,  14'd245,  14'd146,  14'd243,  14'd2422,  14'd934,  14'd448,  14'd755,  -14'd971,  -14'd1924,  -14'd814,  14'd836,  
-14'd175,  14'd420,  -14'd1900,  14'd1397,  -14'd52,  14'd842,  14'd283,  -14'd264,  14'd1009,  14'd1188,  14'd1379,  14'd196,  -14'd721,  -14'd1345,  -14'd694,  14'd393,  
14'd1558,  14'd877,  14'd736,  14'd882,  14'd697,  -14'd448,  14'd336,  -14'd781,  14'd1953,  -14'd189,  14'd553,  14'd1215,  14'd399,  14'd761,  -14'd67,  14'd387,  
14'd1035,  14'd27,  14'd785,  -14'd1621,  -14'd226,  -14'd699,  14'd494,  14'd764,  14'd356,  14'd1336,  -14'd103,  14'd1715,  14'd851,  14'd1800,  14'd362,  -14'd352,  
14'd1081,  14'd65,  -14'd808,  -14'd1108,  -14'd1288,  14'd1010,  14'd371,  -14'd716,  -14'd206,  -14'd745,  -14'd350,  14'd591,  14'd845,  14'd1558,  -14'd180,  -14'd442,  

-14'd2445,  14'd1090,  14'd133,  -14'd1453,  -14'd28,  14'd125,  14'd547,  -14'd1697,  -14'd455,  -14'd1713,  -14'd2137,  14'd384,  -14'd1940,  14'd650,  -14'd997,  14'd848,  
-14'd825,  14'd264,  14'd1724,  14'd76,  14'd817,  -14'd987,  -14'd426,  -14'd965,  -14'd839,  -14'd964,  -14'd1187,  14'd761,  -14'd714,  14'd124,  -14'd942,  -14'd165,  
14'd357,  14'd2143,  -14'd323,  -14'd875,  14'd964,  14'd1053,  -14'd1056,  -14'd1696,  14'd1022,  14'd95,  -14'd359,  14'd518,  -14'd1823,  14'd1854,  -14'd152,  14'd435,  
14'd657,  14'd884,  -14'd610,  14'd127,  -14'd275,  14'd1224,  -14'd58,  -14'd970,  14'd832,  -14'd303,  -14'd378,  -14'd767,  -14'd219,  14'd1284,  -14'd661,  14'd801,  
14'd1451,  14'd1732,  -14'd1858,  -14'd388,  14'd198,  14'd1224,  14'd421,  -14'd589,  14'd115,  -14'd1332,  14'd717,  14'd757,  14'd736,  -14'd641,  -14'd187,  -14'd305,  
14'd256,  14'd269,  14'd1017,  -14'd232,  -14'd195,  -14'd45,  14'd804,  -14'd1366,  -14'd2320,  14'd630,  -14'd374,  14'd1663,  -14'd1316,  14'd893,  14'd1149,  -14'd1177,  
14'd220,  -14'd1237,  14'd462,  -14'd501,  14'd700,  -14'd664,  14'd281,  -14'd42,  14'd1027,  14'd6,  -14'd441,  14'd1707,  -14'd576,  14'd550,  -14'd248,  -14'd1295,  
14'd367,  14'd328,  14'd562,  -14'd550,  14'd781,  -14'd919,  14'd769,  -14'd931,  -14'd797,  14'd362,  -14'd482,  -14'd1167,  14'd1470,  -14'd550,  14'd1378,  -14'd1694,  
-14'd283,  -14'd1627,  14'd578,  -14'd512,  14'd1598,  -14'd401,  14'd241,  14'd648,  -14'd484,  -14'd734,  -14'd2138,  14'd1171,  -14'd1494,  14'd77,  -14'd1141,  14'd405,  
14'd526,  14'd1059,  -14'd827,  -14'd1216,  -14'd1095,  -14'd498,  14'd923,  -14'd756,  14'd764,  -14'd559,  14'd1422,  -14'd1427,  -14'd137,  -14'd599,  -14'd118,  -14'd716,  
14'd204,  -14'd722,  14'd440,  14'd847,  -14'd1502,  14'd169,  14'd237,  14'd557,  14'd574,  14'd888,  -14'd1,  -14'd491,  -14'd757,  14'd1911,  14'd1110,  -14'd900,  
-14'd42,  -14'd254,  14'd540,  14'd1186,  -14'd807,  14'd1543,  14'd322,  -14'd624,  14'd143,  14'd447,  -14'd1201,  14'd593,  14'd1010,  -14'd759,  -14'd259,  14'd536,  
14'd679,  -14'd383,  -14'd986,  14'd1787,  14'd129,  -14'd180,  -14'd381,  14'd770,  -14'd1161,  -14'd764,  14'd1032,  -14'd942,  14'd984,  14'd588,  14'd1429,  14'd883,  
14'd988,  -14'd652,  14'd2071,  14'd398,  -14'd1052,  14'd1794,  14'd855,  14'd619,  14'd135,  -14'd1321,  14'd94,  14'd265,  -14'd51,  -14'd526,  14'd232,  -14'd185,  
-14'd542,  -14'd568,  -14'd1091,  14'd66,  -14'd151,  14'd259,  14'd133,  14'd283,  -14'd1179,  -14'd686,  14'd311,  -14'd495,  14'd1234,  14'd812,  -14'd353,  14'd636,  
14'd1152,  -14'd838,  -14'd554,  14'd813,  14'd1017,  14'd258,  14'd394,  14'd94,  -14'd1195,  14'd622,  14'd862,  -14'd20,  14'd535,  14'd1189,  14'd878,  14'd1127,  
-14'd1711,  14'd790,  14'd120,  14'd173,  14'd1411,  -14'd1084,  14'd770,  -14'd358,  14'd380,  14'd13,  14'd628,  14'd423,  14'd456,  -14'd314,  -14'd1136,  14'd741,  
-14'd265,  14'd96,  -14'd499,  14'd684,  14'd28,  -14'd718,  -14'd225,  14'd277,  -14'd406,  -14'd44,  -14'd858,  -14'd1170,  -14'd151,  -14'd899,  14'd714,  -14'd200,  
-14'd769,  14'd45,  -14'd631,  -14'd249,  -14'd45,  -14'd273,  -14'd378,  14'd1670,  -14'd1752,  -14'd738,  14'd572,  14'd583,  -14'd849,  -14'd1333,  -14'd372,  -14'd751,  
14'd712,  -14'd884,  -14'd2431,  -14'd34,  -14'd1535,  14'd683,  -14'd527,  14'd362,  -14'd814,  -14'd846,  14'd204,  -14'd37,  -14'd336,  -14'd1157,  14'd695,  14'd1176,  
-14'd167,  14'd1220,  14'd1256,  14'd139,  14'd1161,  14'd905,  -14'd275,  14'd1146,  -14'd673,  -14'd1099,  14'd660,  14'd957,  -14'd244,  -14'd847,  14'd100,  14'd77,  
14'd785,  14'd292,  14'd739,  -14'd324,  14'd1330,  -14'd556,  14'd277,  -14'd942,  -14'd81,  -14'd210,  -14'd290,  -14'd356,  14'd9,  14'd626,  -14'd1424,  14'd503,  
-14'd477,  14'd293,  -14'd755,  -14'd1459,  14'd285,  -14'd1260,  -14'd234,  -14'd602,  -14'd1121,  14'd1329,  -14'd517,  -14'd290,  -14'd244,  14'd1344,  14'd404,  -14'd480,  
-14'd493,  14'd337,  14'd1102,  14'd1076,  14'd1328,  -14'd1042,  -14'd199,  -14'd223,  -14'd311,  14'd514,  14'd213,  14'd979,  14'd26,  14'd258,  -14'd468,  -14'd132,  
-14'd775,  -14'd1138,  14'd478,  14'd1688,  14'd454,  14'd427,  14'd635,  -14'd664,  -14'd1163,  14'd1593,  -14'd415,  14'd470,  -14'd513,  -14'd1584,  14'd99,  14'd332,  

14'd17,  -14'd1068,  -14'd290,  14'd603,  -14'd277,  -14'd159,  14'd161,  14'd568,  -14'd333,  -14'd167,  14'd2419,  -14'd1192,  14'd997,  -14'd565,  14'd279,  14'd1452,  
14'd817,  -14'd52,  14'd402,  -14'd162,  -14'd692,  14'd1290,  14'd178,  14'd195,  14'd70,  -14'd1151,  14'd2112,  -14'd42,  -14'd929,  -14'd1245,  -14'd1431,  -14'd673,  
-14'd379,  14'd654,  14'd751,  14'd421,  -14'd298,  -14'd590,  -14'd380,  -14'd661,  -14'd1116,  -14'd1225,  14'd1217,  14'd555,  -14'd143,  -14'd231,  14'd13,  14'd1582,  
14'd2017,  -14'd378,  -14'd1549,  -14'd385,  -14'd371,  -14'd847,  -14'd1024,  14'd1097,  14'd713,  14'd1100,  14'd1030,  -14'd209,  14'd38,  -14'd1604,  -14'd81,  14'd183,  
14'd155,  14'd254,  14'd978,  14'd1478,  -14'd331,  14'd818,  -14'd142,  14'd826,  14'd1178,  14'd852,  14'd43,  -14'd278,  -14'd571,  14'd470,  14'd612,  14'd46,  
-14'd1624,  14'd721,  14'd1629,  14'd519,  14'd7,  -14'd1192,  14'd178,  -14'd477,  -14'd572,  14'd547,  -14'd451,  14'd782,  -14'd2110,  -14'd1198,  14'd1230,  14'd1045,  
-14'd926,  14'd422,  -14'd563,  -14'd841,  -14'd335,  -14'd288,  14'd1660,  -14'd1137,  14'd495,  -14'd318,  14'd1831,  -14'd269,  14'd291,  -14'd553,  -14'd2147,  -14'd141,  
-14'd507,  14'd1999,  14'd77,  14'd82,  14'd209,  14'd531,  14'd1441,  -14'd1199,  -14'd522,  -14'd232,  14'd791,  -14'd789,  14'd338,  14'd1296,  -14'd2050,  14'd3,  
-14'd731,  14'd976,  -14'd641,  -14'd518,  14'd1046,  14'd567,  -14'd1034,  14'd106,  14'd915,  -14'd86,  14'd1596,  -14'd962,  14'd805,  14'd950,  14'd940,  14'd440,  
-14'd1235,  -14'd1339,  -14'd1229,  14'd269,  14'd605,  -14'd404,  14'd619,  -14'd989,  14'd218,  -14'd258,  -14'd958,  -14'd283,  -14'd499,  14'd184,  14'd1552,  -14'd119,  
14'd405,  -14'd856,  14'd637,  -14'd939,  -14'd1184,  14'd1246,  14'd183,  14'd609,  14'd402,  -14'd632,  -14'd1743,  14'd436,  14'd9,  -14'd851,  14'd610,  -14'd471,  
14'd1279,  -14'd80,  -14'd216,  14'd797,  14'd1101,  14'd1225,  -14'd585,  -14'd270,  14'd871,  14'd299,  14'd213,  -14'd211,  14'd163,  -14'd899,  14'd101,  -14'd42,  
14'd831,  -14'd356,  14'd130,  -14'd1382,  -14'd583,  -14'd200,  -14'd876,  -14'd237,  14'd311,  14'd1624,  -14'd812,  -14'd924,  14'd1048,  14'd454,  -14'd1512,  -14'd447,  
14'd1129,  -14'd759,  -14'd89,  -14'd155,  14'd1037,  14'd1341,  14'd280,  -14'd1050,  -14'd278,  -14'd1025,  -14'd133,  14'd531,  -14'd3099,  14'd1180,  -14'd584,  14'd114,  
14'd389,  14'd528,  14'd2636,  -14'd689,  -14'd1617,  14'd83,  14'd1637,  14'd705,  14'd1014,  14'd1205,  -14'd1462,  14'd2279,  -14'd1400,  -14'd365,  -14'd964,  -14'd57,  
14'd1251,  14'd1272,  14'd1302,  -14'd1017,  -14'd1265,  -14'd6,  -14'd349,  14'd1254,  -14'd145,  -14'd391,  -14'd1486,  14'd220,  -14'd349,  -14'd77,  -14'd314,  14'd189,  
-14'd356,  -14'd84,  14'd1339,  14'd550,  -14'd1111,  -14'd1332,  14'd1479,  -14'd507,  14'd529,  -14'd100,  14'd1228,  14'd1257,  14'd594,  14'd306,  -14'd277,  -14'd364,  
-14'd1527,  -14'd713,  14'd1225,  -14'd35,  -14'd993,  -14'd291,  14'd208,  -14'd107,  -14'd249,  14'd651,  14'd533,  14'd218,  -14'd442,  14'd1224,  -14'd161,  14'd78,  
14'd1803,  14'd1168,  -14'd390,  14'd28,  -14'd1357,  -14'd1335,  14'd1055,  14'd28,  14'd605,  14'd685,  14'd537,  14'd1256,  14'd1363,  14'd243,  -14'd377,  14'd200,  
14'd857,  14'd363,  14'd606,  14'd494,  14'd719,  14'd629,  -14'd648,  14'd1109,  14'd1278,  -14'd915,  14'd704,  14'd1601,  14'd222,  14'd902,  14'd814,  14'd1209,  
-14'd983,  14'd690,  14'd260,  -14'd1001,  -14'd2154,  14'd968,  14'd373,  14'd571,  -14'd2080,  -14'd30,  -14'd483,  14'd1004,  -14'd1252,  14'd1386,  -14'd1296,  14'd873,  
14'd779,  14'd1314,  -14'd986,  -14'd727,  -14'd157,  -14'd940,  14'd785,  -14'd254,  14'd1462,  -14'd683,  -14'd715,  14'd22,  14'd646,  14'd1061,  14'd1643,  14'd484,  
-14'd812,  14'd233,  14'd877,  -14'd1508,  -14'd813,  14'd262,  14'd567,  14'd520,  -14'd1028,  -14'd445,  -14'd355,  -14'd875,  14'd815,  -14'd717,  14'd159,  14'd636,  
14'd154,  -14'd605,  14'd1717,  -14'd445,  -14'd998,  -14'd1578,  14'd1136,  -14'd681,  -14'd536,  -14'd587,  14'd406,  -14'd197,  -14'd1200,  14'd1024,  -14'd80,  -14'd775,  
-14'd1521,  -14'd645,  -14'd1847,  -14'd1384,  14'd73,  -14'd151,  -14'd588,  14'd277,  -14'd2389,  -14'd1172,  -14'd1159,  -14'd2159,  -14'd765,  14'd673,  -14'd1307,  -14'd228,  

14'd164,  14'd374,  -14'd361,  14'd42,  14'd475,  14'd143,  -14'd27,  14'd1538,  14'd184,  -14'd1151,  14'd1202,  -14'd90,  -14'd477,  -14'd437,  -14'd1103,  -14'd684,  
14'd356,  14'd575,  14'd21,  14'd265,  14'd170,  14'd550,  14'd830,  14'd31,  -14'd985,  -14'd1951,  -14'd1503,  14'd362,  -14'd197,  14'd1548,  14'd898,  14'd229,  
14'd1209,  14'd596,  -14'd633,  14'd516,  -14'd812,  14'd196,  -14'd385,  -14'd1297,  14'd1559,  -14'd1609,  -14'd594,  14'd895,  -14'd376,  14'd894,  -14'd190,  14'd159,  
-14'd471,  14'd354,  14'd797,  -14'd1754,  14'd442,  -14'd190,  -14'd3,  14'd494,  14'd42,  14'd1595,  14'd226,  -14'd23,  14'd900,  14'd1536,  -14'd1507,  14'd1494,  
14'd194,  14'd668,  14'd353,  14'd411,  14'd318,  14'd462,  14'd1037,  -14'd912,  14'd738,  14'd482,  14'd992,  14'd685,  14'd690,  -14'd1400,  -14'd340,  14'd79,  
14'd143,  -14'd619,  -14'd1965,  14'd1055,  -14'd183,  -14'd114,  14'd306,  -14'd1535,  -14'd7,  -14'd177,  -14'd743,  14'd157,  -14'd721,  -14'd682,  -14'd1466,  -14'd366,  
14'd524,  14'd338,  14'd1605,  14'd34,  -14'd1237,  -14'd703,  -14'd1452,  -14'd40,  -14'd516,  14'd60,  14'd876,  14'd837,  -14'd1163,  14'd390,  14'd362,  14'd718,  
-14'd1178,  -14'd1433,  14'd645,  14'd896,  14'd261,  -14'd327,  -14'd674,  -14'd437,  -14'd475,  -14'd456,  14'd318,  -14'd468,  -14'd1723,  -14'd101,  14'd1322,  -14'd296,  
-14'd1208,  14'd723,  -14'd234,  -14'd405,  -14'd46,  -14'd266,  -14'd338,  14'd86,  14'd346,  -14'd554,  -14'd1058,  14'd477,  -14'd295,  14'd471,  14'd447,  -14'd483,  
14'd360,  14'd1831,  14'd161,  14'd95,  -14'd198,  -14'd810,  -14'd375,  -14'd804,  14'd316,  14'd1236,  -14'd1480,  14'd1266,  14'd315,  -14'd495,  -14'd618,  14'd952,  
14'd959,  14'd1564,  -14'd1214,  14'd228,  -14'd1546,  14'd943,  -14'd391,  -14'd909,  14'd694,  -14'd877,  14'd1298,  -14'd43,  -14'd73,  14'd144,  14'd1407,  -14'd1128,  
14'd450,  14'd1007,  -14'd315,  14'd427,  -14'd284,  -14'd144,  -14'd304,  -14'd406,  14'd1564,  14'd1427,  14'd50,  14'd1254,  14'd1924,  14'd765,  -14'd1571,  14'd111,  
-14'd234,  -14'd365,  -14'd38,  -14'd727,  -14'd622,  -14'd415,  14'd220,  14'd93,  14'd1446,  -14'd134,  14'd177,  14'd833,  14'd763,  14'd9,  -14'd1058,  -14'd542,  
-14'd677,  -14'd811,  14'd447,  14'd646,  -14'd842,  -14'd387,  -14'd688,  14'd120,  -14'd455,  14'd609,  -14'd1095,  14'd544,  14'd609,  14'd1116,  14'd139,  -14'd847,  
14'd1744,  -14'd202,  -14'd1931,  14'd440,  14'd324,  14'd1902,  -14'd1405,  -14'd263,  14'd1316,  -14'd439,  14'd586,  -14'd245,  14'd472,  14'd661,  -14'd568,  14'd333,  
14'd1539,  -14'd254,  14'd1694,  14'd609,  -14'd768,  -14'd660,  14'd237,  -14'd615,  14'd164,  -14'd777,  -14'd834,  14'd104,  14'd832,  14'd958,  -14'd464,  14'd170,  
14'd1627,  14'd1083,  -14'd151,  14'd8,  -14'd588,  -14'd1578,  -14'd67,  14'd111,  14'd1077,  14'd185,  14'd226,  14'd1692,  14'd1239,  14'd475,  -14'd198,  14'd6,  
-14'd187,  14'd309,  -14'd551,  14'd191,  14'd437,  14'd925,  14'd242,  14'd674,  14'd861,  -14'd1416,  14'd462,  -14'd509,  14'd868,  -14'd830,  -14'd856,  14'd575,  
-14'd408,  -14'd114,  -14'd106,  14'd1432,  14'd2094,  14'd991,  14'd598,  14'd384,  -14'd1527,  14'd465,  -14'd324,  -14'd139,  -14'd1037,  -14'd787,  14'd1884,  14'd455,  
-14'd319,  -14'd965,  -14'd820,  14'd451,  -14'd850,  14'd265,  -14'd728,  14'd285,  -14'd354,  14'd2096,  14'd1424,  14'd1314,  14'd912,  14'd1136,  -14'd141,  14'd744,  
-14'd3,  -14'd993,  14'd1431,  14'd370,  -14'd6,  14'd375,  14'd730,  14'd939,  -14'd747,  14'd138,  -14'd490,  -14'd1545,  14'd56,  14'd1467,  14'd1260,  14'd128,  
-14'd473,  -14'd197,  -14'd1016,  -14'd344,  -14'd211,  14'd267,  14'd912,  14'd507,  -14'd602,  -14'd1428,  14'd173,  14'd473,  -14'd94,  -14'd620,  -14'd657,  -14'd702,  
-14'd985,  -14'd360,  14'd78,  14'd578,  14'd715,  -14'd654,  -14'd1404,  -14'd50,  -14'd2338,  -14'd1072,  14'd909,  -14'd208,  -14'd743,  -14'd595,  -14'd872,  14'd296,  
-14'd1935,  14'd234,  -14'd371,  14'd8,  -14'd29,  -14'd300,  -14'd382,  14'd523,  -14'd1401,  14'd402,  -14'd744,  14'd209,  -14'd37,  -14'd783,  14'd128,  -14'd594,  
-14'd1358,  -14'd202,  -14'd1393,  14'd946,  14'd304,  -14'd479,  -14'd528,  14'd814,  14'd753,  14'd1301,  14'd1873,  14'd1179,  14'd168,  14'd192,  14'd16,  14'd1814,  

14'd703,  14'd872,  -14'd495,  -14'd918,  -14'd634,  -14'd489,  14'd211,  -14'd1165,  -14'd960,  14'd3,  -14'd29,  14'd82,  -14'd1059,  -14'd1755,  -14'd1266,  -14'd330,  
14'd1228,  14'd480,  -14'd1207,  14'd840,  -14'd1059,  14'd453,  -14'd1151,  14'd412,  14'd754,  -14'd378,  14'd792,  -14'd1316,  -14'd161,  14'd76,  -14'd22,  -14'd71,  
14'd1384,  -14'd684,  -14'd2153,  14'd1410,  -14'd728,  -14'd663,  -14'd586,  -14'd336,  14'd1540,  14'd653,  -14'd1213,  14'd427,  14'd673,  -14'd2355,  -14'd249,  14'd2053,  
-14'd437,  -14'd905,  14'd409,  -14'd425,  14'd1267,  -14'd398,  -14'd1743,  14'd185,  14'd24,  14'd1297,  -14'd1507,  -14'd214,  14'd246,  14'd451,  14'd770,  14'd773,  
-14'd114,  14'd51,  14'd997,  14'd334,  14'd953,  -14'd236,  -14'd1674,  -14'd35,  -14'd761,  14'd958,  -14'd1825,  -14'd434,  -14'd540,  14'd84,  -14'd909,  -14'd594,  
14'd460,  14'd113,  14'd519,  -14'd259,  14'd115,  14'd498,  -14'd609,  14'd253,  -14'd15,  14'd599,  -14'd463,  14'd979,  -14'd793,  14'd253,  -14'd572,  14'd421,  
-14'd293,  14'd1031,  -14'd1097,  -14'd455,  -14'd437,  -14'd688,  -14'd1217,  14'd1412,  -14'd457,  14'd557,  -14'd1819,  14'd342,  14'd747,  14'd1483,  14'd673,  14'd1192,  
-14'd733,  -14'd1224,  14'd562,  -14'd531,  14'd830,  14'd188,  -14'd717,  14'd410,  14'd147,  14'd1001,  -14'd754,  14'd739,  -14'd223,  -14'd334,  14'd1060,  -14'd546,  
-14'd281,  -14'd440,  14'd429,  14'd106,  -14'd1018,  14'd386,  14'd313,  -14'd789,  -14'd1160,  -14'd1745,  -14'd503,  -14'd707,  14'd752,  14'd378,  14'd344,  -14'd513,  
14'd203,  -14'd456,  14'd155,  14'd1081,  -14'd961,  -14'd318,  14'd355,  -14'd735,  14'd566,  -14'd2131,  -14'd911,  -14'd408,  14'd678,  14'd303,  14'd260,  14'd201,  
14'd722,  14'd239,  -14'd877,  14'd369,  14'd1755,  14'd705,  -14'd657,  -14'd371,  14'd844,  14'd1696,  -14'd197,  14'd667,  14'd1091,  14'd172,  14'd319,  -14'd783,  
-14'd818,  14'd629,  14'd1191,  14'd376,  14'd199,  14'd1239,  -14'd893,  14'd1986,  -14'd812,  14'd708,  14'd341,  -14'd65,  14'd1056,  14'd174,  14'd366,  -14'd257,  
14'd312,  14'd474,  14'd1303,  -14'd6,  14'd508,  14'd117,  14'd1712,  14'd638,  -14'd186,  -14'd770,  14'd10,  -14'd29,  14'd130,  14'd72,  14'd1471,  -14'd1197,  
14'd1865,  14'd157,  14'd1638,  -14'd177,  -14'd481,  14'd1345,  14'd2020,  -14'd470,  -14'd782,  -14'd96,  14'd1077,  -14'd1403,  -14'd789,  14'd1214,  -14'd883,  -14'd233,  
14'd2312,  14'd576,  -14'd2026,  14'd341,  -14'd1549,  14'd773,  14'd16,  14'd487,  -14'd201,  -14'd1773,  -14'd1276,  -14'd738,  14'd1821,  14'd1054,  -14'd277,  14'd1213,  
-14'd1672,  -14'd213,  -14'd1341,  14'd397,  14'd3130,  14'd1171,  -14'd1478,  -14'd674,  14'd152,  -14'd175,  -14'd631,  14'd634,  -14'd261,  -14'd1296,  14'd734,  -14'd415,  
-14'd1137,  14'd663,  14'd839,  14'd551,  14'd1467,  -14'd444,  14'd100,  -14'd2,  -14'd104,  14'd603,  14'd920,  14'd194,  -14'd347,  14'd577,  -14'd1882,  14'd561,  
14'd1371,  -14'd805,  14'd945,  14'd355,  14'd324,  14'd868,  -14'd71,  14'd729,  14'd774,  -14'd257,  -14'd798,  14'd775,  -14'd276,  14'd388,  -14'd1940,  -14'd390,  
-14'd507,  14'd684,  14'd874,  -14'd980,  -14'd132,  -14'd1148,  14'd992,  -14'd658,  -14'd226,  14'd878,  -14'd1158,  -14'd247,  -14'd1188,  14'd1107,  -14'd139,  14'd803,  
-14'd458,  -14'd807,  14'd209,  14'd1105,  -14'd691,  -14'd504,  -14'd1131,  -14'd326,  14'd247,  -14'd243,  -14'd1542,  -14'd1377,  -14'd721,  14'd1804,  -14'd411,  -14'd659,  
-14'd371,  14'd110,  -14'd667,  14'd699,  14'd1429,  -14'd716,  -14'd284,  -14'd591,  14'd900,  -14'd371,  14'd82,  -14'd330,  14'd370,  14'd41,  14'd487,  14'd267,  
-14'd665,  -14'd1292,  -14'd0,  14'd1236,  14'd359,  -14'd285,  14'd1581,  14'd1238,  14'd1751,  14'd568,  14'd1370,  -14'd957,  14'd47,  14'd237,  14'd221,  14'd792,  
-14'd893,  14'd163,  14'd94,  14'd611,  -14'd226,  -14'd80,  -14'd617,  -14'd1242,  -14'd498,  -14'd294,  14'd23,  14'd96,  14'd173,  14'd758,  -14'd637,  14'd883,  
-14'd858,  -14'd1373,  14'd369,  -14'd407,  14'd497,  -14'd84,  14'd591,  14'd897,  14'd606,  14'd302,  -14'd46,  -14'd1138,  14'd150,  14'd800,  14'd904,  14'd1032,  
-14'd353,  -14'd1542,  14'd503,  -14'd45,  -14'd746,  14'd686,  -14'd53,  -14'd1502,  14'd453,  -14'd433,  -14'd646,  14'd1290,  14'd1299,  14'd1362,  14'd902,  14'd223,  

-14'd94,  14'd19,  -14'd1201,  -14'd204,  -14'd15,  -14'd230,  -14'd405,  -14'd96,  -14'd1365,  14'd351,  14'd759,  -14'd792,  -14'd139,  14'd760,  -14'd821,  14'd105,  
14'd251,  14'd170,  -14'd751,  14'd1116,  -14'd503,  -14'd571,  14'd561,  -14'd1044,  14'd1227,  -14'd962,  14'd916,  -14'd1401,  14'd961,  14'd244,  14'd557,  -14'd296,  
-14'd484,  14'd304,  -14'd645,  -14'd1012,  -14'd481,  14'd722,  -14'd1437,  -14'd883,  -14'd1030,  14'd1233,  -14'd1212,  -14'd630,  14'd216,  -14'd144,  -14'd0,  -14'd301,  
-14'd611,  -14'd561,  -14'd389,  -14'd449,  -14'd201,  -14'd442,  -14'd729,  -14'd389,  -14'd650,  14'd851,  14'd907,  -14'd656,  -14'd174,  -14'd9,  14'd67,  14'd536,  
14'd28,  -14'd1084,  -14'd48,  14'd689,  14'd854,  14'd514,  -14'd474,  14'd640,  14'd779,  14'd352,  14'd1043,  -14'd591,  14'd729,  -14'd961,  -14'd98,  14'd744,  
14'd486,  -14'd180,  -14'd94,  14'd743,  -14'd820,  -14'd1305,  -14'd468,  -14'd562,  14'd608,  14'd1461,  14'd403,  14'd488,  14'd51,  -14'd139,  14'd1276,  -14'd345,  
-14'd352,  -14'd142,  -14'd601,  -14'd500,  -14'd98,  -14'd1492,  -14'd91,  14'd452,  -14'd61,  14'd341,  -14'd253,  -14'd607,  14'd579,  -14'd355,  -14'd635,  -14'd579,  
-14'd837,  14'd1334,  -14'd200,  14'd259,  14'd856,  14'd269,  14'd291,  14'd132,  -14'd763,  14'd60,  -14'd154,  -14'd739,  -14'd546,  -14'd752,  -14'd201,  -14'd815,  
14'd1111,  -14'd97,  14'd1115,  14'd406,  14'd427,  -14'd1134,  -14'd872,  -14'd173,  14'd547,  -14'd817,  -14'd208,  -14'd1117,  14'd384,  14'd967,  -14'd458,  -14'd1183,  
14'd470,  14'd722,  14'd84,  14'd970,  -14'd65,  -14'd554,  -14'd1051,  -14'd757,  -14'd1462,  14'd363,  -14'd991,  -14'd691,  -14'd827,  14'd627,  -14'd335,  14'd745,  
14'd1072,  -14'd1709,  14'd677,  -14'd1355,  -14'd472,  14'd830,  14'd327,  -14'd970,  -14'd531,  14'd368,  -14'd198,  -14'd718,  14'd886,  -14'd534,  -14'd489,  -14'd750,  
14'd1428,  -14'd33,  -14'd259,  -14'd401,  -14'd405,  -14'd541,  14'd966,  -14'd207,  -14'd332,  -14'd498,  -14'd710,  -14'd103,  14'd342,  14'd425,  14'd569,  -14'd1619,  
14'd1047,  14'd581,  14'd207,  -14'd1515,  14'd263,  14'd259,  -14'd1687,  14'd140,  14'd140,  14'd1191,  14'd791,  -14'd131,  14'd128,  14'd78,  14'd37,  14'd772,  
-14'd518,  14'd1167,  -14'd1334,  -14'd7,  -14'd861,  -14'd149,  -14'd624,  14'd543,  -14'd477,  14'd524,  14'd1044,  -14'd1036,  -14'd290,  -14'd400,  -14'd61,  14'd715,  
-14'd767,  -14'd142,  -14'd1068,  -14'd1601,  -14'd602,  14'd861,  -14'd377,  -14'd324,  14'd516,  -14'd144,  14'd459,  -14'd595,  -14'd387,  14'd189,  -14'd560,  -14'd1171,  
-14'd615,  14'd216,  14'd184,  -14'd904,  14'd385,  -14'd1017,  14'd1331,  14'd670,  -14'd1080,  14'd297,  14'd90,  14'd749,  -14'd297,  14'd38,  -14'd176,  -14'd488,  
14'd1271,  14'd547,  14'd227,  -14'd909,  -14'd672,  -14'd430,  14'd816,  -14'd1201,  14'd734,  -14'd35,  -14'd441,  -14'd652,  -14'd487,  -14'd1150,  14'd142,  -14'd907,  
-14'd447,  -14'd347,  -14'd1017,  14'd1365,  -14'd124,  14'd1502,  -14'd495,  -14'd743,  -14'd1288,  14'd96,  -14'd1269,  -14'd768,  -14'd739,  -14'd546,  -14'd712,  -14'd718,  
-14'd392,  14'd486,  14'd492,  14'd40,  -14'd250,  -14'd1341,  14'd125,  14'd1152,  14'd361,  -14'd634,  -14'd224,  14'd25,  14'd349,  -14'd273,  14'd361,  14'd774,  
-14'd1069,  -14'd637,  14'd1037,  14'd255,  -14'd28,  -14'd309,  -14'd588,  -14'd572,  -14'd1287,  14'd619,  14'd534,  14'd709,  14'd1240,  -14'd109,  -14'd905,  14'd417,  
-14'd239,  -14'd914,  14'd888,  14'd1089,  -14'd381,  -14'd68,  -14'd1692,  14'd997,  -14'd680,  -14'd737,  -14'd1233,  -14'd836,  -14'd124,  -14'd816,  -14'd638,  -14'd770,  
-14'd43,  -14'd1038,  -14'd93,  14'd16,  -14'd1320,  -14'd312,  -14'd1340,  -14'd182,  -14'd60,  -14'd543,  14'd1245,  -14'd551,  -14'd1307,  14'd190,  -14'd555,  -14'd571,  
-14'd1209,  -14'd517,  14'd37,  14'd106,  14'd85,  -14'd909,  -14'd94,  -14'd1253,  -14'd986,  14'd474,  -14'd861,  14'd966,  14'd70,  -14'd587,  14'd1159,  -14'd1075,  
14'd162,  14'd65,  -14'd229,  14'd1002,  -14'd370,  14'd414,  -14'd618,  14'd613,  -14'd415,  -14'd591,  -14'd289,  -14'd730,  14'd436,  -14'd1619,  -14'd134,  -14'd1387,  
14'd1075,  -14'd553,  -14'd900,  -14'd1391,  -14'd510,  14'd785,  -14'd270,  -14'd106,  -14'd474,  -14'd430,  14'd274,  14'd388,  14'd977,  -14'd1078,  14'd708,  14'd587,  

-14'd277,  14'd185,  14'd1009,  14'd298,  -14'd819,  -14'd749,  14'd649,  14'd1254,  14'd280,  14'd239,  -14'd16,  -14'd427,  14'd879,  14'd1074,  -14'd4,  14'd377,  
-14'd576,  14'd178,  14'd2652,  -14'd1994,  14'd1138,  -14'd1305,  14'd1070,  14'd25,  -14'd731,  14'd132,  -14'd2609,  14'd317,  -14'd11,  14'd2062,  -14'd194,  14'd231,  
14'd465,  14'd315,  14'd1,  -14'd1509,  14'd76,  -14'd969,  14'd2303,  14'd342,  -14'd701,  14'd22,  -14'd828,  -14'd343,  -14'd1288,  14'd2708,  -14'd1002,  -14'd1471,  
-14'd887,  14'd762,  14'd733,  -14'd593,  14'd935,  -14'd473,  14'd1418,  -14'd996,  14'd328,  -14'd361,  14'd239,  -14'd643,  -14'd1503,  14'd1402,  14'd1096,  -14'd1147,  
14'd1164,  14'd1015,  -14'd979,  -14'd374,  14'd33,  14'd2202,  14'd456,  14'd259,  14'd765,  14'd352,  14'd235,  -14'd510,  14'd486,  -14'd440,  -14'd259,  14'd448,  
14'd38,  -14'd464,  14'd72,  14'd594,  14'd540,  14'd181,  14'd441,  -14'd184,  -14'd1237,  -14'd616,  -14'd720,  14'd886,  14'd158,  14'd729,  14'd162,  -14'd627,  
14'd1278,  -14'd1414,  14'd444,  14'd518,  -14'd545,  -14'd1456,  14'd1093,  -14'd43,  -14'd205,  -14'd683,  -14'd1041,  14'd599,  -14'd1405,  14'd2012,  -14'd1189,  -14'd1721,  
14'd79,  14'd1023,  14'd1177,  -14'd327,  -14'd947,  -14'd641,  14'd787,  -14'd610,  14'd601,  14'd83,  -14'd373,  -14'd196,  -14'd742,  14'd1570,  14'd543,  -14'd1914,  
14'd769,  -14'd189,  -14'd525,  -14'd1654,  14'd1103,  -14'd925,  -14'd359,  -14'd239,  -14'd454,  -14'd1917,  -14'd471,  14'd513,  14'd480,  14'd696,  -14'd1468,  -14'd126,  
14'd1410,  14'd275,  14'd379,  -14'd957,  14'd104,  14'd1144,  14'd341,  -14'd626,  14'd1781,  14'd166,  14'd645,  -14'd452,  -14'd626,  -14'd220,  -14'd510,  -14'd651,  
-14'd719,  -14'd669,  -14'd1814,  14'd410,  -14'd1005,  14'd123,  14'd446,  -14'd800,  -14'd247,  -14'd626,  14'd1990,  14'd445,  14'd1428,  14'd635,  14'd439,  -14'd767,  
14'd365,  14'd142,  14'd130,  14'd274,  -14'd1635,  14'd251,  14'd969,  -14'd987,  -14'd168,  14'd1070,  -14'd437,  -14'd799,  14'd1314,  14'd423,  14'd419,  14'd1322,  
-14'd681,  14'd296,  14'd334,  14'd1250,  14'd987,  14'd37,  14'd44,  -14'd144,  -14'd422,  -14'd616,  14'd1075,  -14'd379,  14'd1253,  -14'd642,  -14'd41,  -14'd380,  
-14'd639,  -14'd1659,  14'd621,  14'd412,  14'd837,  14'd822,  14'd511,  14'd494,  14'd1307,  -14'd939,  14'd85,  -14'd343,  -14'd544,  -14'd1535,  -14'd148,  14'd554,  
-14'd859,  -14'd99,  -14'd1061,  14'd1011,  -14'd240,  14'd240,  -14'd133,  -14'd1085,  -14'd1320,  14'd1010,  14'd212,  -14'd282,  14'd824,  -14'd1032,  -14'd110,  14'd522,  
-14'd945,  14'd150,  14'd748,  -14'd1106,  -14'd889,  -14'd591,  -14'd1025,  -14'd39,  14'd724,  -14'd327,  14'd209,  14'd231,  14'd1781,  -14'd37,  14'd843,  -14'd547,  
14'd235,  -14'd450,  -14'd82,  -14'd201,  14'd238,  14'd91,  14'd815,  14'd1040,  -14'd605,  14'd430,  14'd1372,  14'd1344,  -14'd221,  14'd640,  -14'd574,  14'd331,  
14'd766,  -14'd1256,  -14'd1275,  14'd1286,  14'd122,  14'd1645,  -14'd365,  -14'd228,  -14'd1317,  -14'd747,  14'd480,  14'd289,  14'd94,  14'd590,  14'd679,  -14'd162,  
-14'd33,  14'd100,  14'd825,  14'd1404,  -14'd596,  14'd144,  14'd178,  14'd1726,  14'd536,  14'd1081,  14'd1029,  14'd707,  -14'd733,  -14'd151,  14'd1062,  14'd803,  
14'd23,  14'd372,  -14'd844,  14'd444,  14'd184,  -14'd838,  -14'd856,  -14'd594,  -14'd261,  -14'd649,  14'd1050,  -14'd269,  14'd867,  14'd213,  14'd760,  14'd848,  
-14'd112,  -14'd504,  14'd701,  -14'd306,  -14'd652,  -14'd243,  -14'd121,  -14'd4,  -14'd1016,  14'd666,  -14'd1850,  -14'd994,  14'd319,  14'd155,  14'd951,  -14'd583,  
-14'd539,  14'd34,  14'd493,  -14'd426,  -14'd782,  -14'd834,  14'd756,  14'd145,  14'd262,  14'd387,  14'd206,  14'd328,  -14'd1591,  14'd715,  -14'd461,  -14'd433,  
14'd1209,  14'd1899,  -14'd123,  -14'd196,  14'd882,  -14'd376,  -14'd728,  -14'd670,  -14'd2128,  14'd168,  14'd134,  -14'd211,  -14'd1562,  14'd682,  -14'd879,  -14'd743,  
-14'd1160,  14'd1684,  14'd1104,  14'd994,  14'd1491,  14'd79,  -14'd483,  -14'd229,  14'd1110,  14'd1957,  -14'd439,  -14'd1126,  14'd79,  -14'd337,  14'd1465,  -14'd507,  
14'd39,  -14'd461,  -14'd869,  14'd454,  14'd1184,  14'd597,  14'd412,  14'd1115,  -14'd254,  14'd1487,  14'd777,  14'd196,  -14'd1096,  14'd170,  14'd712,  14'd1475,  

-14'd2017,  -14'd34,  14'd157,  14'd297,  14'd361,  14'd613,  14'd84,  -14'd501,  14'd551,  14'd534,  14'd1497,  -14'd1418,  -14'd164,  -14'd457,  14'd2211,  -14'd231,  
-14'd1111,  -14'd1163,  -14'd1522,  -14'd534,  14'd530,  -14'd764,  -14'd900,  14'd1165,  14'd693,  14'd100,  14'd571,  -14'd515,  14'd363,  14'd362,  14'd25,  14'd411,  
14'd213,  -14'd2611,  14'd1140,  14'd1182,  14'd1101,  -14'd1098,  14'd111,  14'd700,  -14'd442,  -14'd239,  14'd390,  14'd987,  -14'd533,  -14'd1227,  14'd1020,  -14'd1251,  
14'd222,  -14'd1486,  14'd444,  14'd570,  -14'd933,  14'd817,  14'd660,  -14'd185,  14'd734,  -14'd255,  14'd562,  14'd412,  -14'd796,  -14'd53,  -14'd424,  -14'd734,  
-14'd1685,  -14'd987,  14'd859,  -14'd520,  -14'd857,  14'd244,  -14'd322,  14'd1130,  -14'd745,  14'd914,  -14'd812,  -14'd737,  -14'd181,  -14'd241,  -14'd365,  -14'd1307,  
14'd290,  14'd723,  14'd285,  -14'd873,  -14'd703,  -14'd717,  -14'd1750,  14'd568,  -14'd1325,  14'd568,  14'd318,  14'd1135,  -14'd919,  14'd846,  -14'd1161,  -14'd1527,  
-14'd763,  -14'd706,  -14'd1866,  -14'd931,  14'd767,  14'd606,  14'd682,  -14'd1830,  -14'd696,  -14'd696,  14'd617,  14'd329,  -14'd648,  -14'd684,  14'd288,  -14'd574,  
-14'd7,  14'd183,  14'd28,  14'd905,  -14'd56,  14'd1044,  -14'd1401,  14'd341,  -14'd1368,  14'd74,  -14'd119,  14'd998,  -14'd355,  -14'd131,  -14'd767,  14'd1595,  
-14'd1135,  14'd522,  -14'd632,  14'd2010,  14'd1061,  14'd1191,  14'd1426,  -14'd795,  -14'd795,  -14'd2,  14'd587,  -14'd477,  -14'd37,  14'd2270,  14'd544,  14'd702,  
-14'd1646,  -14'd2451,  -14'd313,  -14'd1413,  14'd510,  -14'd902,  14'd693,  14'd791,  -14'd948,  14'd408,  -14'd486,  -14'd1464,  -14'd1364,  14'd925,  -14'd874,  14'd216,  
14'd423,  14'd1107,  14'd729,  14'd159,  -14'd407,  -14'd405,  -14'd15,  14'd1063,  -14'd464,  -14'd1422,  14'd1462,  14'd384,  -14'd1553,  14'd1041,  -14'd1221,  -14'd961,  
14'd367,  -14'd16,  -14'd1653,  -14'd1426,  14'd307,  -14'd1121,  14'd1436,  -14'd452,  -14'd678,  14'd879,  -14'd65,  14'd1286,  14'd191,  14'd487,  14'd1208,  14'd1276,  
14'd614,  14'd769,  14'd825,  14'd1403,  -14'd421,  14'd537,  14'd286,  14'd708,  -14'd167,  14'd724,  14'd518,  14'd1234,  14'd1144,  14'd305,  14'd174,  -14'd75,  
14'd210,  -14'd527,  14'd922,  14'd313,  14'd66,  14'd999,  14'd981,  -14'd775,  -14'd43,  -14'd2522,  14'd150,  14'd725,  -14'd1025,  -14'd367,  14'd1275,  -14'd82,  
-14'd1476,  -14'd1392,  14'd1880,  14'd846,  14'd323,  14'd521,  14'd57,  -14'd802,  -14'd1493,  -14'd140,  -14'd296,  14'd985,  -14'd569,  -14'd253,  -14'd944,  -14'd804,  
-14'd400,  14'd562,  14'd1073,  -14'd1638,  -14'd1439,  14'd387,  14'd1372,  -14'd496,  -14'd733,  -14'd123,  14'd674,  14'd265,  -14'd630,  14'd571,  -14'd358,  14'd858,  
-14'd49,  14'd429,  -14'd391,  -14'd948,  14'd12,  -14'd494,  14'd1531,  -14'd497,  14'd582,  -14'd758,  14'd378,  14'd122,  14'd741,  -14'd501,  14'd446,  14'd125,  
14'd353,  14'd114,  14'd972,  14'd738,  -14'd976,  -14'd178,  14'd326,  14'd1479,  14'd73,  -14'd721,  14'd350,  -14'd363,  14'd23,  14'd255,  -14'd413,  14'd111,  
14'd605,  14'd467,  14'd1098,  -14'd100,  -14'd962,  -14'd276,  14'd1315,  14'd1270,  14'd1190,  -14'd2363,  14'd1841,  -14'd361,  14'd1249,  -14'd1808,  -14'd765,  -14'd262,  
14'd1176,  14'd478,  -14'd499,  -14'd748,  -14'd595,  -14'd56,  -14'd408,  14'd1216,  -14'd1816,  -14'd2820,  -14'd72,  14'd129,  14'd854,  14'd1185,  14'd1805,  14'd889,  
-14'd282,  -14'd1583,  -14'd1282,  -14'd1384,  -14'd868,  -14'd1743,  14'd1731,  14'd230,  -14'd1057,  14'd924,  14'd277,  -14'd820,  -14'd559,  14'd134,  14'd206,  -14'd118,  
-14'd530,  14'd312,  14'd1017,  -14'd239,  -14'd157,  14'd1042,  14'd2481,  14'd1053,  14'd535,  14'd1133,  -14'd451,  14'd389,  14'd570,  14'd1049,  -14'd711,  -14'd486,  
-14'd694,  14'd1070,  14'd1901,  -14'd1988,  14'd1350,  -14'd2553,  14'd493,  14'd764,  14'd1223,  -14'd220,  -14'd824,  -14'd1735,  -14'd997,  14'd526,  14'd1364,  -14'd1020,  
14'd180,  -14'd764,  -14'd784,  -14'd380,  -14'd887,  -14'd1902,  -14'd46,  14'd415,  -14'd603,  -14'd1683,  -14'd1443,  -14'd2150,  -14'd2030,  -14'd159,  -14'd1378,  -14'd372,  
-14'd695,  -14'd587,  14'd987,  -14'd1017,  -14'd1951,  -14'd793,  -14'd35,  14'd539,  -14'd791,  -14'd1128,  -14'd1080,  -14'd1339,  -14'd1256,  -14'd1248,  -14'd822,  -14'd1554,  

-14'd508,  -14'd932,  14'd381,  14'd202,  14'd134,  -14'd155,  -14'd1644,  14'd1674,  14'd133,  14'd1069,  -14'd442,  -14'd726,  -14'd320,  -14'd237,  14'd1807,  14'd1569,  
-14'd520,  -14'd1309,  14'd372,  14'd868,  14'd179,  14'd405,  -14'd1606,  14'd560,  -14'd899,  14'd1428,  14'd1564,  14'd216,  14'd1347,  -14'd960,  14'd878,  14'd321,  
14'd850,  -14'd21,  -14'd341,  14'd536,  14'd198,  14'd254,  14'd123,  -14'd660,  -14'd1624,  14'd104,  14'd818,  14'd159,  14'd665,  -14'd3680,  -14'd1395,  14'd1108,  
14'd1549,  -14'd44,  -14'd312,  14'd218,  -14'd315,  14'd1426,  14'd832,  -14'd251,  14'd1326,  -14'd733,  14'd674,  14'd870,  -14'd407,  -14'd1421,  -14'd418,  -14'd169,  
14'd1085,  -14'd1416,  14'd1496,  -14'd295,  -14'd2,  -14'd406,  14'd645,  -14'd588,  14'd382,  14'd556,  -14'd590,  -14'd57,  -14'd1175,  -14'd327,  -14'd942,  14'd447,  
-14'd512,  14'd649,  -14'd286,  -14'd196,  14'd1147,  14'd865,  -14'd1048,  14'd742,  14'd1183,  -14'd370,  14'd459,  14'd735,  14'd1410,  14'd23,  14'd60,  -14'd1081,  
-14'd1062,  -14'd901,  -14'd1768,  14'd1430,  14'd408,  -14'd778,  -14'd1651,  -14'd550,  -14'd1231,  -14'd371,  14'd580,  14'd833,  14'd1325,  -14'd532,  14'd461,  -14'd576,  
14'd1050,  -14'd674,  -14'd1388,  14'd1269,  14'd1038,  14'd401,  -14'd1436,  14'd1145,  -14'd638,  14'd308,  14'd214,  14'd137,  14'd435,  -14'd431,  14'd351,  14'd1041,  
14'd745,  14'd336,  -14'd1407,  14'd401,  14'd645,  14'd211,  14'd1468,  14'd1470,  14'd886,  14'd793,  14'd1781,  -14'd734,  14'd629,  14'd90,  -14'd144,  14'd554,  
14'd182,  -14'd2237,  -14'd640,  14'd364,  -14'd1050,  14'd423,  -14'd1082,  14'd1130,  14'd803,  14'd1102,  14'd322,  -14'd381,  14'd1078,  -14'd128,  -14'd363,  -14'd505,  
-14'd1054,  14'd1282,  -14'd448,  14'd979,  14'd1107,  -14'd703,  14'd214,  14'd458,  14'd2501,  14'd539,  14'd1266,  14'd400,  -14'd54,  14'd930,  -14'd5,  14'd86,  
-14'd875,  -14'd200,  -14'd468,  14'd589,  14'd48,  -14'd1804,  -14'd1749,  -14'd785,  -14'd1420,  -14'd243,  14'd1110,  -14'd97,  14'd1320,  -14'd449,  -14'd86,  14'd805,  
-14'd15,  -14'd647,  14'd1245,  14'd308,  -14'd1587,  14'd1412,  14'd925,  14'd220,  -14'd928,  14'd1893,  14'd629,  14'd859,  14'd612,  -14'd1452,  -14'd702,  14'd1327,  
14'd439,  14'd687,  -14'd1353,  14'd2,  14'd728,  14'd1551,  -14'd348,  14'd1210,  -14'd366,  -14'd649,  -14'd297,  14'd603,  14'd150,  14'd192,  14'd552,  14'd306,  
-14'd1330,  -14'd563,  -14'd828,  -14'd32,  14'd1405,  -14'd676,  -14'd641,  -14'd108,  14'd300,  -14'd196,  14'd1087,  14'd455,  14'd1460,  14'd53,  14'd795,  -14'd1227,  
-14'd299,  14'd306,  -14'd1153,  -14'd1381,  14'd525,  -14'd202,  -14'd729,  14'd261,  14'd1109,  -14'd39,  14'd640,  14'd384,  -14'd381,  -14'd1084,  -14'd1790,  -14'd803,  
-14'd2001,  -14'd1381,  14'd700,  14'd580,  -14'd819,  -14'd942,  -14'd480,  -14'd1479,  14'd146,  14'd679,  -14'd14,  14'd158,  -14'd991,  -14'd1433,  14'd211,  14'd1561,  
-14'd1495,  14'd263,  -14'd66,  14'd246,  14'd321,  -14'd422,  14'd151,  -14'd811,  14'd1774,  -14'd4,  14'd226,  14'd244,  14'd530,  -14'd1828,  -14'd450,  -14'd582,  
-14'd273,  14'd721,  14'd686,  -14'd1414,  -14'd1139,  14'd888,  -14'd101,  -14'd480,  -14'd460,  14'd762,  14'd45,  14'd307,  -14'd5,  -14'd1193,  -14'd1294,  -14'd391,  
14'd895,  -14'd576,  -14'd671,  14'd384,  -14'd216,  -14'd406,  -14'd887,  14'd2007,  -14'd845,  14'd633,  -14'd260,  14'd169,  14'd890,  14'd658,  -14'd295,  14'd518,  
14'd736,  14'd1131,  -14'd753,  -14'd427,  14'd1483,  14'd858,  14'd1251,  -14'd1786,  14'd952,  14'd1004,  -14'd227,  14'd127,  14'd329,  -14'd905,  -14'd1203,  14'd298,  
-14'd400,  -14'd666,  14'd331,  -14'd1430,  -14'd412,  14'd1049,  14'd1171,  -14'd250,  14'd849,  14'd1671,  -14'd767,  -14'd884,  -14'd449,  14'd992,  -14'd475,  14'd807,  
14'd126,  14'd1646,  14'd867,  -14'd166,  -14'd556,  14'd57,  14'd1837,  -14'd374,  14'd489,  14'd1131,  -14'd436,  -14'd848,  14'd436,  -14'd708,  14'd763,  14'd20,  
14'd94,  -14'd1243,  14'd126,  -14'd692,  14'd411,  14'd159,  14'd91,  -14'd273,  14'd803,  -14'd694,  -14'd1274,  -14'd2131,  -14'd2231,  14'd1140,  14'd146,  14'd474,  
14'd490,  -14'd538,  14'd1069,  -14'd1192,  -14'd422,  -14'd652,  -14'd769,  -14'd885,  14'd634,  -14'd836,  -14'd301,  -14'd435,  14'd409,  -14'd1249,  -14'd1123,  14'd76,  

14'd1591,  14'd171,  14'd140,  -14'd59,  -14'd461,  -14'd966,  14'd771,  14'd35,  14'd422,  -14'd465,  -14'd550,  -14'd589,  14'd23,  14'd149,  -14'd1893,  -14'd817,  
14'd2241,  14'd310,  14'd1084,  -14'd257,  -14'd38,  14'd613,  14'd1294,  -14'd66,  14'd206,  -14'd106,  14'd863,  14'd530,  14'd80,  14'd403,  -14'd495,  14'd1606,  
14'd1914,  14'd110,  14'd148,  14'd1235,  -14'd323,  -14'd1184,  14'd371,  14'd556,  -14'd396,  -14'd250,  14'd820,  14'd90,  14'd1516,  -14'd910,  14'd304,  14'd366,  
-14'd871,  14'd841,  14'd1581,  14'd316,  -14'd136,  14'd994,  -14'd2451,  -14'd868,  -14'd1635,  -14'd410,  -14'd577,  -14'd1012,  14'd754,  -14'd560,  14'd179,  -14'd545,  
14'd453,  -14'd413,  14'd201,  -14'd48,  14'd1673,  -14'd1251,  -14'd438,  -14'd1102,  -14'd2136,  -14'd767,  -14'd250,  -14'd1117,  14'd1322,  14'd384,  14'd21,  14'd2532,  
14'd1293,  -14'd1690,  14'd1519,  -14'd254,  -14'd52,  14'd1409,  -14'd312,  14'd998,  -14'd41,  -14'd170,  -14'd1247,  -14'd852,  14'd68,  14'd548,  14'd205,  -14'd1033,  
-14'd214,  -14'd1014,  -14'd135,  -14'd546,  -14'd276,  -14'd103,  -14'd335,  -14'd471,  -14'd873,  14'd40,  14'd381,  14'd1237,  -14'd1001,  -14'd674,  -14'd28,  -14'd635,  
-14'd295,  14'd452,  -14'd833,  -14'd904,  14'd1282,  14'd766,  14'd66,  14'd350,  14'd1007,  14'd1801,  14'd1149,  -14'd133,  -14'd352,  -14'd619,  -14'd273,  14'd322,  
-14'd381,  -14'd80,  -14'd288,  -14'd379,  14'd485,  -14'd1089,  -14'd1857,  14'd376,  -14'd841,  14'd2069,  14'd1071,  -14'd323,  14'd223,  -14'd1325,  -14'd1085,  14'd795,  
-14'd577,  -14'd199,  -14'd619,  -14'd564,  14'd1862,  14'd951,  -14'd888,  14'd676,  -14'd373,  14'd581,  14'd373,  14'd183,  -14'd91,  14'd189,  -14'd753,  14'd768,  
14'd211,  14'd36,  14'd178,  -14'd531,  14'd857,  -14'd13,  -14'd907,  -14'd439,  -14'd1117,  14'd577,  -14'd1279,  14'd431,  -14'd1257,  14'd365,  14'd1412,  -14'd430,  
-14'd675,  14'd260,  -14'd549,  14'd230,  14'd1016,  14'd966,  -14'd681,  -14'd912,  14'd221,  14'd285,  14'd65,  14'd60,  -14'd723,  -14'd1116,  14'd148,  -14'd187,  
14'd300,  -14'd828,  14'd302,  14'd1327,  14'd918,  14'd106,  -14'd96,  14'd1279,  14'd1914,  -14'd188,  -14'd207,  14'd440,  -14'd1937,  -14'd453,  -14'd354,  14'd46,  
14'd1425,  -14'd636,  -14'd633,  -14'd372,  -14'd548,  14'd393,  -14'd663,  -14'd185,  14'd902,  14'd2576,  14'd179,  -14'd607,  14'd937,  14'd436,  -14'd2113,  14'd267,  
14'd611,  14'd598,  -14'd1209,  -14'd442,  14'd1588,  14'd671,  -14'd339,  -14'd967,  14'd486,  14'd1613,  14'd652,  14'd938,  -14'd799,  -14'd5,  -14'd853,  -14'd240,  
14'd993,  14'd470,  -14'd419,  14'd1072,  -14'd126,  -14'd1367,  14'd424,  -14'd252,  -14'd972,  14'd877,  -14'd1462,  14'd598,  14'd75,  14'd748,  14'd405,  14'd510,  
14'd1597,  14'd1477,  14'd558,  14'd1661,  -14'd44,  -14'd318,  14'd72,  -14'd608,  14'd1400,  14'd1431,  -14'd126,  14'd1085,  -14'd477,  14'd680,  14'd467,  -14'd1235,  
14'd1036,  14'd1276,  -14'd71,  14'd397,  14'd1397,  14'd237,  -14'd1182,  -14'd358,  -14'd692,  -14'd467,  14'd975,  14'd346,  -14'd551,  14'd852,  -14'd217,  14'd833,  
-14'd779,  14'd849,  -14'd1026,  -14'd347,  14'd621,  -14'd1503,  -14'd985,  14'd217,  -14'd951,  -14'd375,  -14'd221,  -14'd162,  14'd230,  -14'd345,  14'd2010,  -14'd713,  
14'd17,  -14'd450,  14'd731,  -14'd178,  -14'd1669,  14'd1362,  -14'd1376,  14'd1185,  14'd491,  14'd86,  -14'd51,  14'd1050,  14'd1119,  14'd827,  -14'd112,  14'd289,  
14'd1232,  14'd70,  14'd301,  14'd735,  -14'd1238,  14'd769,  14'd1,  14'd1232,  14'd930,  14'd1230,  -14'd29,  14'd694,  14'd29,  14'd2373,  -14'd44,  -14'd475,  
14'd331,  14'd226,  14'd142,  14'd1172,  14'd904,  14'd90,  -14'd781,  14'd960,  14'd224,  -14'd413,  14'd811,  -14'd611,  14'd679,  14'd857,  14'd2016,  -14'd198,  
-14'd667,  -14'd434,  -14'd1374,  14'd51,  14'd1002,  14'd599,  -14'd680,  14'd251,  -14'd571,  -14'd1373,  -14'd223,  -14'd193,  14'd920,  -14'd2654,  14'd523,  -14'd106,  
14'd610,  14'd234,  14'd354,  -14'd231,  14'd324,  14'd1296,  14'd70,  14'd1761,  14'd199,  -14'd329,  -14'd420,  14'd1290,  14'd671,  14'd197,  -14'd76,  14'd562,  
14'd332,  14'd871,  14'd1249,  -14'd2,  -14'd807,  14'd308,  14'd958,  14'd677,  14'd1383,  14'd454,  -14'd1130,  14'd2205,  -14'd859,  -14'd446,  14'd11,  14'd8,  

-14'd988,  14'd810,  -14'd645,  14'd462,  14'd1787,  -14'd239,  -14'd1427,  14'd793,  -14'd1014,  14'd325,  -14'd200,  14'd230,  -14'd167,  14'd884,  -14'd230,  14'd2060,  
-14'd1127,  14'd807,  14'd333,  14'd1009,  14'd662,  14'd891,  -14'd694,  -14'd187,  14'd493,  14'd998,  -14'd1394,  14'd771,  -14'd338,  -14'd1565,  14'd1854,  14'd2394,  
-14'd953,  -14'd140,  14'd1116,  14'd516,  -14'd289,  -14'd917,  14'd186,  14'd573,  14'd63,  14'd72,  -14'd1009,  14'd353,  14'd729,  14'd868,  -14'd1223,  14'd1214,  
-14'd507,  -14'd1693,  14'd127,  -14'd19,  14'd178,  -14'd497,  14'd1414,  -14'd807,  -14'd23,  -14'd649,  14'd564,  14'd1187,  -14'd1152,  14'd2727,  14'd137,  -14'd1704,  
-14'd1488,  14'd622,  14'd1096,  -14'd1128,  -14'd1150,  -14'd490,  14'd337,  -14'd1238,  14'd279,  -14'd331,  -14'd1501,  -14'd1125,  -14'd1621,  14'd1217,  -14'd1500,  -14'd1107,  
14'd992,  14'd1237,  -14'd834,  -14'd664,  14'd689,  -14'd328,  -14'd506,  14'd678,  -14'd331,  -14'd1140,  14'd351,  14'd49,  14'd393,  -14'd1119,  14'd814,  14'd1115,  
14'd147,  14'd480,  -14'd785,  -14'd911,  14'd288,  14'd670,  -14'd427,  -14'd612,  14'd166,  14'd2047,  14'd797,  14'd1174,  -14'd331,  14'd30,  14'd1075,  14'd377,  
14'd1898,  14'd566,  14'd1934,  14'd705,  -14'd1074,  -14'd754,  14'd91,  -14'd49,  14'd189,  14'd559,  -14'd272,  14'd1288,  14'd153,  -14'd897,  14'd172,  14'd23,  
14'd1548,  -14'd793,  14'd638,  14'd1357,  14'd62,  14'd1517,  14'd1782,  -14'd238,  -14'd1052,  14'd792,  14'd334,  14'd548,  14'd159,  14'd2944,  -14'd545,  -14'd530,  
14'd915,  -14'd311,  14'd269,  14'd420,  14'd1225,  14'd1456,  14'd215,  -14'd1663,  -14'd3,  -14'd1126,  14'd401,  -14'd532,  14'd478,  14'd1767,  -14'd1815,  -14'd1326,  
-14'd2188,  -14'd450,  -14'd1035,  14'd32,  14'd24,  -14'd968,  14'd799,  14'd398,  14'd1364,  14'd520,  -14'd272,  -14'd793,  -14'd490,  -14'd655,  -14'd1773,  14'd571,  
14'd670,  14'd126,  -14'd30,  14'd51,  -14'd365,  -14'd278,  -14'd1327,  14'd1269,  -14'd965,  14'd6,  -14'd357,  -14'd705,  14'd751,  14'd1498,  14'd630,  14'd22,  
14'd705,  -14'd844,  -14'd974,  -14'd192,  14'd114,  -14'd354,  -14'd203,  14'd1150,  -14'd2749,  14'd425,  14'd898,  -14'd355,  14'd1406,  -14'd346,  14'd768,  -14'd983,  
-14'd3,  -14'd602,  14'd897,  14'd1539,  14'd401,  14'd677,  -14'd266,  14'd790,  -14'd467,  14'd471,  14'd1275,  14'd463,  14'd791,  -14'd567,  -14'd940,  14'd188,  
-14'd598,  -14'd1578,  -14'd111,  -14'd1419,  14'd997,  14'd249,  -14'd125,  14'd502,  -14'd137,  14'd375,  14'd534,  14'd401,  14'd1473,  14'd127,  -14'd1092,  -14'd203,  
-14'd2379,  -14'd1998,  14'd367,  14'd840,  14'd833,  -14'd3,  -14'd1519,  14'd1179,  14'd1185,  -14'd115,  14'd51,  -14'd2072,  -14'd711,  -14'd206,  -14'd445,  -14'd980,  
-14'd1185,  14'd182,  14'd663,  -14'd508,  14'd416,  14'd279,  -14'd742,  -14'd1084,  -14'd295,  14'd636,  14'd391,  -14'd959,  -14'd595,  -14'd1416,  -14'd90,  -14'd290,  
-14'd958,  14'd899,  14'd288,  -14'd648,  -14'd1052,  -14'd620,  -14'd297,  14'd795,  14'd319,  14'd859,  14'd957,  14'd164,  -14'd1344,  -14'd522,  14'd184,  14'd223,  
-14'd779,  -14'd237,  -14'd74,  -14'd1337,  -14'd637,  14'd905,  -14'd727,  14'd335,  14'd428,  -14'd875,  14'd972,  -14'd607,  -14'd91,  14'd1282,  -14'd733,  14'd185,  
14'd197,  14'd1093,  14'd94,  -14'd1096,  14'd409,  14'd96,  14'd200,  -14'd667,  -14'd270,  -14'd612,  14'd8,  -14'd820,  14'd950,  14'd93,  14'd231,  14'd446,  
-14'd1218,  -14'd1251,  -14'd325,  -14'd74,  14'd306,  -14'd337,  14'd2030,  -14'd892,  -14'd86,  -14'd45,  -14'd645,  14'd1077,  14'd1530,  -14'd810,  14'd850,  -14'd426,  
14'd1888,  -14'd285,  14'd529,  -14'd550,  14'd1238,  14'd229,  14'd1007,  -14'd1130,  14'd636,  -14'd214,  -14'd73,  14'd1013,  -14'd717,  -14'd33,  14'd791,  14'd811,  
14'd794,  14'd1606,  14'd580,  14'd48,  14'd233,  14'd399,  14'd191,  14'd234,  -14'd432,  -14'd842,  -14'd84,  14'd861,  14'd102,  14'd584,  -14'd948,  14'd312,  
-14'd491,  -14'd525,  14'd397,  -14'd783,  -14'd541,  -14'd1329,  14'd1176,  14'd108,  -14'd915,  14'd403,  14'd645,  14'd369,  -14'd146,  14'd969,  -14'd433,  14'd147,  
14'd769,  14'd857,  14'd894,  14'd846,  14'd738,  -14'd1802,  14'd1526,  -14'd589,  -14'd242,  14'd510,  14'd149,  14'd641,  -14'd656,  14'd750,  -14'd619,  -14'd749,  

-14'd211,  -14'd237,  -14'd515,  -14'd375,  -14'd1216,  14'd379,  -14'd1748,  -14'd75,  -14'd1919,  -14'd663,  14'd1960,  -14'd761,  -14'd9,  -14'd1361,  14'd494,  14'd513,  
-14'd25,  14'd563,  -14'd1738,  14'd727,  14'd1457,  14'd1197,  -14'd790,  14'd1223,  14'd1359,  -14'd214,  -14'd223,  14'd1226,  14'd594,  -14'd1422,  14'd591,  -14'd364,  
-14'd249,  14'd961,  14'd822,  -14'd286,  14'd666,  14'd820,  -14'd1667,  14'd628,  14'd857,  -14'd1220,  -14'd753,  14'd981,  14'd595,  -14'd1815,  14'd534,  14'd607,  
14'd792,  -14'd312,  14'd1584,  14'd148,  -14'd486,  14'd276,  14'd1121,  14'd1156,  14'd452,  14'd1589,  14'd663,  -14'd242,  14'd1945,  -14'd970,  14'd474,  14'd188,  
-14'd489,  -14'd2777,  -14'd458,  14'd159,  -14'd422,  14'd1108,  14'd765,  -14'd458,  -14'd400,  14'd1253,  14'd969,  -14'd1016,  -14'd589,  -14'd899,  14'd85,  -14'd438,  
-14'd682,  -14'd1207,  14'd22,  -14'd992,  14'd86,  -14'd337,  14'd254,  -14'd1349,  -14'd699,  -14'd1539,  14'd559,  -14'd865,  -14'd680,  14'd59,  -14'd829,  14'd359,  
14'd25,  14'd145,  -14'd1707,  14'd196,  -14'd93,  14'd942,  14'd551,  -14'd908,  -14'd433,  14'd843,  -14'd241,  -14'd536,  14'd109,  -14'd169,  -14'd1845,  14'd1212,  
-14'd1170,  14'd1857,  -14'd693,  -14'd1136,  -14'd242,  14'd156,  14'd260,  -14'd479,  14'd179,  14'd688,  14'd389,  -14'd818,  14'd261,  14'd1941,  -14'd935,  -14'd443,  
14'd457,  14'd742,  14'd219,  -14'd245,  14'd46,  14'd1671,  14'd1462,  -14'd418,  14'd999,  -14'd670,  -14'd718,  14'd1141,  -14'd71,  14'd2471,  14'd1056,  14'd93,  
-14'd2422,  14'd1839,  14'd1354,  14'd376,  14'd444,  -14'd281,  -14'd802,  -14'd989,  -14'd163,  -14'd1654,  14'd434,  -14'd1670,  -14'd2170,  14'd753,  14'd2224,  -14'd934,  
-14'd1254,  -14'd972,  -14'd1011,  -14'd222,  -14'd982,  -14'd1764,  14'd1120,  -14'd1038,  -14'd755,  14'd632,  14'd302,  14'd288,  -14'd1075,  -14'd1010,  14'd194,  -14'd778,  
-14'd105,  14'd100,  -14'd973,  14'd59,  -14'd83,  14'd246,  14'd626,  -14'd996,  14'd1512,  -14'd111,  -14'd1111,  14'd880,  14'd487,  -14'd3040,  -14'd307,  14'd373,  
-14'd325,  14'd221,  -14'd654,  -14'd1445,  -14'd15,  -14'd1290,  14'd920,  -14'd378,  14'd322,  14'd953,  -14'd102,  -14'd749,  -14'd232,  14'd692,  -14'd141,  -14'd61,  
14'd741,  14'd328,  14'd682,  14'd1330,  -14'd642,  14'd344,  14'd342,  -14'd259,  14'd70,  -14'd1937,  -14'd682,  14'd1567,  -14'd566,  14'd229,  14'd547,  -14'd1954,  
14'd1880,  -14'd160,  -14'd369,  14'd1344,  -14'd1793,  14'd481,  -14'd353,  -14'd26,  -14'd196,  -14'd337,  -14'd91,  14'd1057,  -14'd163,  14'd288,  14'd904,  -14'd1602,  
14'd1127,  -14'd1090,  14'd962,  14'd915,  -14'd2761,  14'd83,  14'd1474,  -14'd13,  14'd708,  14'd322,  14'd1048,  14'd37,  -14'd543,  -14'd167,  -14'd102,  14'd598,  
14'd83,  -14'd1715,  -14'd128,  -14'd360,  -14'd1379,  -14'd305,  -14'd898,  -14'd18,  14'd486,  14'd622,  -14'd563,  14'd1556,  14'd1392,  -14'd575,  -14'd559,  14'd17,  
14'd1110,  -14'd915,  14'd614,  -14'd216,  -14'd702,  14'd1144,  -14'd616,  14'd869,  -14'd274,  -14'd495,  -14'd1897,  14'd452,  14'd1006,  14'd606,  14'd828,  -14'd210,  
14'd574,  14'd110,  14'd483,  14'd1046,  -14'd163,  14'd686,  14'd749,  14'd1192,  14'd1688,  14'd1393,  -14'd591,  14'd110,  -14'd92,  -14'd1096,  -14'd711,  -14'd545,  
14'd1107,  14'd736,  -14'd1766,  14'd573,  -14'd61,  14'd724,  14'd155,  14'd756,  -14'd37,  14'd908,  14'd1317,  14'd148,  14'd530,  14'd513,  14'd462,  14'd369,  
14'd330,  -14'd722,  14'd1329,  -14'd943,  -14'd724,  14'd553,  -14'd21,  14'd153,  -14'd746,  -14'd144,  14'd319,  -14'd321,  -14'd182,  14'd824,  -14'd324,  14'd1067,  
-14'd554,  14'd657,  -14'd1402,  -14'd407,  -14'd162,  14'd1063,  14'd849,  -14'd18,  14'd921,  -14'd1361,  14'd1031,  -14'd1000,  14'd418,  14'd363,  14'd809,  14'd288,  
-14'd502,  14'd1113,  14'd550,  -14'd376,  -14'd587,  -14'd724,  -14'd782,  14'd535,  -14'd989,  -14'd904,  14'd285,  -14'd876,  14'd717,  14'd1222,  -14'd632,  -14'd805,  
-14'd1632,  14'd601,  -14'd25,  14'd708,  -14'd161,  14'd460,  -14'd333,  14'd471,  -14'd838,  -14'd205,  -14'd44,  -14'd1100,  14'd99,  14'd379,  14'd243,  14'd235,  
-14'd275,  -14'd691,  -14'd2037,  -14'd707,  -14'd431,  14'd487,  14'd600,  14'd299,  -14'd2323,  14'd3358,  14'd641,  14'd301,  -14'd640,  -14'd449,  -14'd705,  14'd1132,  

-14'd738,  -14'd507,  14'd628,  -14'd937,  -14'd138,  -14'd728,  14'd3290,  -14'd928,  14'd1209,  14'd400,  14'd596,  14'd149,  -14'd143,  14'd564,  14'd1203,  14'd1622,  
-14'd1382,  14'd473,  14'd796,  -14'd1419,  -14'd1889,  14'd520,  14'd2912,  14'd120,  -14'd1345,  14'd89,  14'd711,  14'd783,  14'd1111,  14'd1729,  -14'd629,  -14'd202,  
14'd654,  -14'd453,  14'd1035,  -14'd1835,  -14'd223,  -14'd702,  14'd1821,  -14'd43,  -14'd1448,  -14'd1807,  14'd626,  14'd1099,  -14'd1736,  14'd1911,  -14'd564,  -14'd2856,  
14'd2976,  14'd533,  -14'd1581,  -14'd1010,  -14'd342,  14'd84,  14'd1453,  -14'd518,  -14'd1038,  -14'd1184,  -14'd50,  14'd345,  14'd179,  14'd1029,  -14'd1566,  -14'd1240,  
14'd821,  14'd1403,  -14'd467,  -14'd102,  -14'd1754,  -14'd481,  14'd113,  -14'd708,  14'd402,  14'd59,  -14'd527,  -14'd698,  -14'd1481,  -14'd49,  14'd205,  14'd292,  
14'd1023,  -14'd670,  14'd1016,  -14'd62,  14'd167,  -14'd1376,  14'd2534,  -14'd1166,  -14'd385,  14'd767,  14'd1750,  -14'd738,  14'd160,  -14'd737,  14'd453,  14'd1135,  
-14'd1025,  14'd583,  14'd97,  -14'd245,  14'd1046,  -14'd601,  14'd1370,  -14'd1473,  -14'd893,  -14'd715,  14'd1241,  14'd155,  14'd368,  -14'd464,  -14'd2197,  -14'd363,  
14'd1959,  14'd1154,  14'd897,  -14'd1057,  -14'd1671,  14'd1,  -14'd1071,  -14'd399,  -14'd324,  14'd490,  -14'd806,  14'd56,  14'd1045,  14'd469,  14'd344,  14'd136,  
14'd1616,  14'd1846,  -14'd582,  14'd666,  -14'd354,  14'd1384,  -14'd839,  -14'd849,  14'd1102,  14'd856,  14'd286,  14'd552,  14'd349,  14'd537,  14'd139,  14'd95,  
-14'd19,  -14'd1292,  14'd414,  14'd930,  14'd757,  -14'd1674,  -14'd309,  -14'd135,  -14'd7,  -14'd31,  14'd146,  14'd1305,  14'd1044,  -14'd1321,  14'd924,  14'd345,  
14'd219,  -14'd1466,  -14'd28,  -14'd263,  -14'd431,  -14'd972,  14'd2811,  -14'd433,  -14'd508,  -14'd793,  14'd296,  14'd1269,  -14'd2076,  -14'd2211,  14'd938,  -14'd1321,  
14'd1455,  -14'd1421,  -14'd1039,  -14'd627,  -14'd556,  14'd1113,  -14'd1128,  -14'd423,  14'd967,  -14'd1384,  14'd396,  14'd203,  -14'd1045,  -14'd161,  -14'd183,  14'd167,  
14'd1520,  14'd564,  -14'd54,  -14'd435,  -14'd241,  -14'd928,  -14'd12,  -14'd202,  -14'd246,  -14'd223,  -14'd1954,  -14'd588,  14'd713,  -14'd1186,  -14'd378,  -14'd576,  
-14'd32,  14'd1002,  -14'd803,  -14'd826,  -14'd176,  14'd1345,  14'd325,  -14'd983,  14'd645,  14'd1230,  -14'd328,  14'd513,  -14'd111,  14'd78,  -14'd202,  -14'd363,  
-14'd576,  -14'd182,  14'd706,  14'd1428,  -14'd637,  14'd286,  -14'd93,  -14'd124,  -14'd725,  14'd482,  -14'd1530,  14'd792,  14'd746,  -14'd58,  14'd888,  14'd0,  
14'd478,  14'd295,  14'd545,  14'd224,  14'd742,  14'd533,  14'd1355,  14'd972,  -14'd118,  14'd277,  -14'd873,  14'd589,  -14'd190,  14'd238,  -14'd147,  14'd22,  
14'd24,  -14'd725,  14'd325,  14'd1316,  14'd160,  -14'd681,  14'd240,  -14'd1378,  14'd354,  14'd136,  14'd672,  -14'd607,  14'd413,  14'd840,  -14'd41,  14'd536,  
14'd679,  -14'd1003,  14'd83,  14'd568,  -14'd1764,  -14'd568,  -14'd1040,  14'd1390,  14'd928,  14'd1381,  -14'd739,  -14'd690,  14'd1567,  -14'd983,  14'd212,  -14'd7,  
14'd1556,  -14'd1153,  -14'd1191,  14'd339,  -14'd1483,  -14'd439,  -14'd996,  14'd732,  -14'd648,  -14'd386,  14'd1432,  14'd190,  14'd1887,  14'd903,  14'd446,  -14'd1410,  
14'd238,  -14'd173,  14'd847,  14'd578,  -14'd54,  -14'd707,  14'd613,  14'd788,  14'd370,  14'd1070,  -14'd788,  -14'd69,  14'd1996,  -14'd398,  -14'd195,  14'd777,  
-14'd597,  14'd675,  14'd15,  14'd1786,  14'd626,  14'd1385,  -14'd971,  14'd380,  14'd1263,  14'd503,  14'd702,  -14'd1657,  -14'd289,  -14'd827,  -14'd272,  14'd495,  
14'd156,  -14'd820,  14'd29,  14'd391,  -14'd402,  -14'd1372,  14'd1102,  -14'd623,  14'd489,  14'd915,  14'd144,  -14'd1301,  14'd946,  -14'd880,  -14'd748,  14'd198,  
-14'd591,  14'd129,  -14'd866,  14'd26,  -14'd963,  14'd506,  -14'd69,  -14'd536,  -14'd161,  14'd1777,  -14'd362,  14'd123,  14'd982,  -14'd1352,  14'd409,  14'd1408,  
-14'd2337,  -14'd782,  -14'd818,  14'd363,  14'd196,  14'd1075,  -14'd703,  -14'd1471,  -14'd645,  14'd1112,  -14'd782,  -14'd981,  -14'd685,  -14'd675,  -14'd1626,  14'd883,  
-14'd577,  -14'd96,  -14'd371,  -14'd377,  14'd443,  -14'd1048,  -14'd1673,  14'd268,  -14'd418,  -14'd614,  14'd952,  -14'd1231,  14'd156,  -14'd123,  -14'd283,  -14'd173,  

-14'd500,  -14'd1837,  -14'd135,  14'd701,  14'd802,  -14'd165,  -14'd1433,  14'd362,  -14'd312,  14'd232,  14'd798,  -14'd191,  -14'd338,  -14'd666,  -14'd472,  -14'd1858,  
-14'd222,  -14'd724,  -14'd1650,  14'd1337,  -14'd385,  14'd861,  -14'd690,  14'd1570,  14'd226,  14'd1224,  -14'd5,  -14'd555,  -14'd661,  -14'd946,  14'd1202,  -14'd1071,  
-14'd467,  -14'd116,  14'd266,  14'd1522,  -14'd1008,  14'd442,  -14'd732,  -14'd271,  -14'd276,  14'd400,  -14'd798,  -14'd221,  14'd1007,  14'd604,  14'd1284,  14'd1034,  
14'd23,  -14'd530,  14'd1228,  14'd141,  -14'd269,  -14'd485,  -14'd11,  14'd1262,  -14'd120,  14'd1440,  14'd428,  -14'd1342,  -14'd715,  -14'd2657,  14'd1222,  14'd1347,  
14'd464,  14'd463,  14'd1521,  -14'd112,  14'd239,  14'd766,  -14'd1392,  14'd1173,  14'd529,  -14'd326,  -14'd1471,  14'd768,  14'd805,  14'd607,  14'd1286,  -14'd1346,  
-14'd865,  -14'd736,  14'd10,  -14'd374,  14'd1399,  14'd461,  -14'd1151,  -14'd22,  14'd131,  14'd571,  -14'd879,  -14'd812,  14'd1403,  14'd802,  -14'd1649,  14'd643,  
14'd1043,  14'd1137,  14'd1307,  -14'd79,  -14'd575,  14'd1815,  -14'd381,  14'd123,  -14'd448,  14'd767,  14'd1831,  -14'd1139,  14'd254,  14'd406,  14'd613,  14'd192,  
-14'd1688,  14'd1937,  14'd348,  -14'd5,  14'd164,  14'd1342,  14'd5,  -14'd582,  14'd289,  -14'd305,  -14'd688,  -14'd1239,  -14'd971,  14'd906,  14'd1165,  14'd683,  
-14'd2208,  14'd1950,  14'd1259,  14'd1348,  14'd1456,  14'd886,  -14'd2002,  14'd944,  -14'd33,  -14'd396,  14'd187,  -14'd1159,  -14'd613,  -14'd767,  14'd656,  14'd332,  
14'd844,  14'd1260,  14'd1185,  14'd749,  -14'd735,  14'd1752,  14'd1096,  14'd460,  -14'd122,  -14'd415,  -14'd34,  -14'd264,  -14'd556,  14'd115,  14'd1285,  14'd798,  
-14'd1004,  -14'd634,  14'd361,  -14'd1512,  -14'd505,  -14'd809,  -14'd1507,  -14'd627,  -14'd263,  -14'd109,  -14'd814,  14'd418,  -14'd45,  -14'd510,  -14'd676,  -14'd305,  
14'd727,  -14'd768,  14'd318,  -14'd623,  14'd468,  14'd766,  14'd284,  -14'd137,  -14'd161,  -14'd481,  14'd994,  -14'd100,  -14'd1001,  14'd1263,  14'd916,  14'd999,  
14'd112,  14'd31,  -14'd366,  -14'd201,  14'd941,  14'd547,  14'd738,  14'd1088,  -14'd470,  -14'd936,  -14'd606,  -14'd492,  -14'd293,  14'd232,  -14'd302,  -14'd459,  
-14'd152,  14'd1301,  14'd351,  14'd366,  -14'd19,  -14'd431,  14'd195,  -14'd617,  14'd966,  -14'd6,  14'd508,  -14'd429,  -14'd455,  14'd943,  14'd1750,  -14'd971,  
14'd2689,  14'd1327,  14'd745,  -14'd550,  14'd464,  -14'd1447,  -14'd593,  -14'd729,  -14'd257,  -14'd640,  -14'd1684,  -14'd100,  14'd687,  -14'd225,  14'd493,  -14'd160,  
14'd1551,  -14'd33,  14'd465,  14'd317,  14'd1123,  -14'd730,  14'd307,  -14'd1430,  14'd1181,  14'd418,  -14'd665,  14'd890,  -14'd1682,  14'd400,  -14'd147,  14'd54,  
14'd1767,  -14'd775,  14'd57,  -14'd126,  -14'd1347,  14'd580,  14'd2066,  -14'd595,  14'd1183,  -14'd41,  14'd652,  14'd1337,  14'd539,  14'd548,  -14'd710,  -14'd220,  
-14'd89,  -14'd1277,  -14'd704,  -14'd51,  14'd1355,  14'd874,  -14'd68,  -14'd325,  14'd235,  14'd1043,  14'd1109,  14'd24,  14'd676,  14'd1717,  -14'd147,  -14'd12,  
-14'd867,  14'd124,  -14'd1301,  14'd794,  14'd141,  -14'd1653,  -14'd1518,  -14'd655,  -14'd183,  14'd121,  -14'd1338,  14'd541,  -14'd454,  -14'd994,  -14'd652,  -14'd1588,  
14'd68,  -14'd147,  14'd1429,  -14'd749,  14'd198,  -14'd834,  -14'd1139,  -14'd723,  -14'd1112,  -14'd699,  14'd773,  -14'd130,  -14'd5,  -14'd1839,  -14'd384,  14'd300,  
-14'd90,  14'd150,  14'd424,  -14'd270,  14'd167,  14'd1250,  -14'd1316,  14'd1250,  -14'd160,  -14'd62,  14'd250,  14'd239,  14'd451,  14'd1111,  14'd137,  -14'd347,  
-14'd694,  14'd933,  14'd754,  14'd229,  -14'd340,  14'd402,  -14'd220,  -14'd163,  14'd539,  -14'd1054,  14'd396,  14'd89,  -14'd219,  14'd1579,  14'd1330,  14'd517,  
14'd511,  -14'd1199,  14'd1061,  -14'd475,  14'd909,  14'd86,  -14'd1101,  -14'd23,  -14'd665,  -14'd284,  14'd129,  -14'd65,  14'd261,  -14'd1160,  14'd1419,  14'd447,  
-14'd597,  -14'd924,  -14'd577,  -14'd117,  14'd251,  14'd444,  14'd211,  14'd471,  -14'd504,  -14'd1570,  14'd1536,  14'd868,  14'd1107,  14'd500,  -14'd948,  -14'd111,  
14'd1325,  -14'd357,  14'd768,  -14'd1378,  -14'd1274,  -14'd499,  14'd380,  14'd211,  14'd420,  -14'd1682,  -14'd261,  14'd564,  -14'd939,  -14'd136,  -14'd1642,  -14'd982,  

14'd165,  -14'd205,  14'd1867,  -14'd373,  14'd156,  -14'd668,  14'd1412,  -14'd922,  14'd979,  14'd473,  -14'd341,  -14'd616,  -14'd724,  14'd1112,  -14'd559,  -14'd1754,  
-14'd126,  -14'd894,  14'd39,  14'd550,  14'd241,  14'd690,  14'd2748,  14'd97,  14'd84,  -14'd1135,  14'd213,  14'd373,  14'd372,  14'd148,  -14'd779,  -14'd1136,  
14'd543,  14'd1501,  -14'd814,  -14'd123,  14'd338,  -14'd428,  -14'd295,  -14'd160,  14'd1264,  -14'd993,  14'd809,  -14'd464,  14'd1283,  -14'd251,  -14'd1767,  -14'd895,  
14'd484,  14'd1680,  -14'd851,  14'd989,  -14'd829,  14'd1501,  -14'd494,  -14'd649,  -14'd285,  -14'd992,  14'd80,  14'd839,  14'd1388,  -14'd462,  14'd505,  14'd1175,  
14'd1150,  14'd1663,  -14'd123,  14'd742,  -14'd262,  -14'd747,  -14'd606,  14'd750,  -14'd1469,  -14'd277,  -14'd336,  -14'd774,  14'd2818,  14'd314,  14'd427,  14'd1151,  
14'd1033,  -14'd409,  14'd1400,  14'd1016,  -14'd631,  14'd100,  -14'd292,  14'd193,  14'd1810,  14'd1885,  -14'd1389,  14'd130,  14'd2423,  14'd885,  14'd1661,  -14'd346,  
-14'd760,  14'd726,  14'd647,  -14'd345,  14'd244,  -14'd803,  -14'd1234,  -14'd484,  14'd21,  14'd305,  -14'd35,  -14'd151,  -14'd1011,  -14'd14,  14'd1322,  14'd83,  
14'd188,  -14'd138,  -14'd508,  -14'd1098,  -14'd842,  -14'd1074,  -14'd617,  -14'd971,  14'd953,  14'd995,  14'd2107,  -14'd775,  14'd10,  -14'd648,  -14'd159,  14'd406,  
-14'd1395,  14'd115,  -14'd614,  -14'd534,  -14'd1144,  14'd1,  -14'd412,  -14'd2369,  -14'd556,  14'd529,  -14'd399,  14'd84,  14'd1075,  -14'd1295,  -14'd948,  14'd566,  
14'd849,  -14'd1112,  -14'd1278,  -14'd548,  14'd660,  14'd840,  -14'd1339,  14'd544,  -14'd701,  14'd1889,  14'd358,  14'd662,  14'd652,  -14'd491,  14'd499,  14'd132,  
-14'd593,  14'd1465,  14'd1104,  14'd1539,  14'd573,  14'd492,  -14'd2742,  -14'd858,  14'd8,  14'd473,  -14'd969,  -14'd264,  14'd149,  14'd1933,  14'd1233,  14'd188,  
-14'd409,  14'd790,  14'd6,  14'd635,  -14'd629,  -14'd146,  14'd275,  -14'd165,  -14'd815,  -14'd519,  14'd522,  14'd741,  -14'd468,  14'd1201,  14'd203,  -14'd26,  
-14'd1838,  -14'd1308,  -14'd1295,  -14'd26,  14'd848,  14'd935,  14'd558,  -14'd234,  14'd949,  -14'd2401,  -14'd317,  14'd1047,  -14'd169,  -14'd1434,  -14'd193,  -14'd1086,  
-14'd920,  14'd1007,  -14'd1535,  14'd618,  14'd1611,  -14'd1583,  -14'd395,  14'd59,  14'd676,  14'd881,  14'd164,  14'd252,  14'd152,  14'd480,  -14'd610,  -14'd64,  
-14'd1160,  -14'd1176,  -14'd771,  14'd608,  14'd848,  14'd1269,  -14'd2183,  -14'd80,  14'd196,  14'd2308,  14'd413,  14'd928,  14'd896,  14'd202,  -14'd20,  -14'd762,  
-14'd241,  -14'd253,  14'd1253,  -14'd297,  14'd660,  14'd124,  14'd677,  14'd597,  -14'd455,  -14'd561,  -14'd835,  14'd413,  -14'd448,  14'd591,  -14'd413,  -14'd616,  
14'd1167,  14'd108,  14'd1138,  -14'd144,  -14'd349,  -14'd717,  -14'd919,  14'd1241,  14'd478,  14'd1046,  -14'd390,  14'd1610,  -14'd325,  14'd1439,  14'd1167,  14'd250,  
-14'd599,  14'd311,  -14'd1000,  -14'd324,  14'd1254,  14'd1158,  14'd12,  14'd612,  -14'd830,  -14'd617,  14'd113,  14'd1033,  -14'd1092,  -14'd2664,  14'd792,  14'd1065,  
-14'd1101,  -14'd372,  -14'd1014,  -14'd1434,  14'd1436,  -14'd72,  -14'd866,  -14'd1730,  14'd334,  -14'd326,  14'd893,  -14'd1171,  14'd316,  14'd638,  14'd1325,  14'd1156,  
-14'd712,  -14'd918,  14'd2311,  -14'd388,  -14'd500,  -14'd226,  -14'd188,  -14'd1124,  14'd634,  -14'd950,  -14'd11,  14'd360,  -14'd40,  14'd63,  -14'd1653,  -14'd768,  
14'd1008,  -14'd1214,  -14'd2,  -14'd1082,  14'd166,  14'd539,  -14'd103,  14'd869,  14'd1735,  -14'd898,  -14'd929,  14'd34,  14'd76,  14'd1568,  -14'd13,  14'd35,  
14'd1320,  14'd510,  14'd249,  14'd729,  14'd698,  -14'd1278,  -14'd1318,  -14'd350,  -14'd211,  -14'd304,  -14'd356,  -14'd7,  14'd938,  -14'd13,  14'd1401,  14'd510,  
-14'd79,  -14'd158,  -14'd1094,  -14'd294,  -14'd453,  14'd622,  14'd504,  14'd375,  -14'd621,  -14'd2281,  -14'd44,  14'd27,  14'd599,  -14'd1751,  14'd759,  14'd75,  
-14'd814,  -14'd989,  -14'd1301,  -14'd1441,  -14'd716,  14'd249,  -14'd521,  14'd1052,  14'd1046,  -14'd1896,  14'd875,  14'd716,  14'd839,  14'd1200,  -14'd516,  -14'd326,  
-14'd121,  14'd517,  -14'd2139,  -14'd244,  -14'd1043,  14'd222,  14'd453,  14'd988,  -14'd379,  -14'd3706,  14'd115,  -14'd63,  -14'd544,  -14'd843,  -14'd241,  -14'd662,  

-14'd552,  14'd329,  14'd1095,  -14'd313,  -14'd300,  14'd449,  14'd1561,  -14'd303,  14'd639,  14'd1000,  -14'd968,  14'd637,  14'd930,  14'd2352,  -14'd522,  14'd274,  
14'd766,  14'd446,  14'd1043,  -14'd463,  -14'd611,  14'd1033,  14'd1342,  14'd707,  14'd416,  14'd226,  14'd616,  14'd884,  14'd1386,  14'd698,  -14'd829,  14'd1353,  
14'd8,  14'd414,  -14'd161,  14'd79,  -14'd369,  14'd153,  14'd661,  14'd823,  14'd824,  -14'd7,  -14'd370,  14'd578,  14'd375,  -14'd449,  14'd655,  14'd375,  
-14'd673,  -14'd310,  14'd82,  -14'd58,  14'd808,  -14'd560,  -14'd734,  -14'd130,  -14'd1373,  -14'd982,  -14'd224,  -14'd1305,  -14'd508,  -14'd1296,  -14'd667,  -14'd773,  
-14'd1116,  14'd2252,  14'd674,  14'd2,  -14'd310,  14'd853,  14'd139,  14'd88,  -14'd1263,  -14'd1237,  14'd190,  14'd1257,  -14'd566,  14'd1687,  14'd358,  14'd2046,  
-14'd734,  14'd690,  14'd450,  -14'd953,  14'd854,  14'd148,  -14'd512,  -14'd82,  14'd500,  14'd859,  -14'd804,  14'd61,  14'd1739,  14'd955,  -14'd1359,  -14'd272,  
14'd852,  -14'd496,  -14'd131,  -14'd208,  14'd1328,  14'd130,  -14'd1049,  -14'd440,  -14'd1424,  14'd474,  -14'd437,  14'd256,  -14'd124,  14'd951,  -14'd186,  -14'd436,  
-14'd1313,  14'd89,  14'd45,  -14'd357,  14'd243,  -14'd760,  -14'd558,  14'd354,  14'd311,  -14'd683,  14'd958,  14'd514,  -14'd748,  14'd1097,  -14'd342,  14'd377,  
-14'd1385,  -14'd626,  14'd481,  -14'd685,  -14'd25,  -14'd453,  -14'd132,  14'd1490,  14'd727,  14'd489,  14'd278,  -14'd1351,  -14'd397,  -14'd1203,  14'd792,  -14'd427,  
-14'd1016,  14'd584,  14'd235,  -14'd375,  14'd312,  14'd39,  -14'd665,  14'd26,  14'd545,  14'd2110,  14'd394,  14'd800,  14'd417,  -14'd632,  14'd681,  14'd1398,  
14'd81,  14'd472,  -14'd1355,  -14'd641,  14'd691,  14'd934,  14'd962,  14'd644,  -14'd1119,  14'd1054,  -14'd751,  14'd952,  -14'd1870,  -14'd983,  14'd680,  14'd346,  
-14'd232,  14'd178,  14'd1443,  -14'd180,  14'd666,  14'd346,  -14'd1321,  -14'd1325,  14'd124,  14'd753,  14'd230,  14'd1336,  -14'd358,  -14'd650,  -14'd1534,  14'd416,  
-14'd1487,  14'd1799,  14'd82,  14'd549,  14'd1308,  14'd201,  14'd151,  14'd1119,  14'd84,  14'd1511,  14'd1058,  14'd89,  -14'd522,  -14'd1013,  -14'd793,  14'd361,  
-14'd1444,  14'd583,  -14'd380,  -14'd104,  14'd43,  14'd836,  -14'd1237,  -14'd2,  14'd339,  14'd994,  -14'd95,  -14'd524,  -14'd333,  -14'd722,  -14'd426,  14'd96,  
14'd415,  -14'd952,  -14'd86,  14'd924,  14'd414,  14'd91,  14'd90,  -14'd20,  14'd1280,  -14'd514,  14'd231,  14'd3,  -14'd740,  14'd474,  -14'd1248,  14'd1677,  
14'd1130,  14'd913,  14'd120,  14'd261,  -14'd669,  14'd894,  14'd1265,  14'd1282,  14'd465,  -14'd776,  14'd886,  14'd1129,  14'd1123,  14'd1665,  14'd708,  14'd1344,  
14'd653,  14'd953,  14'd591,  14'd109,  14'd336,  14'd944,  14'd533,  -14'd1616,  14'd693,  14'd1524,  -14'd240,  14'd452,  -14'd303,  14'd121,  14'd835,  14'd418,  
-14'd361,  14'd858,  -14'd1481,  14'd352,  14'd530,  14'd628,  14'd193,  14'd3,  -14'd724,  -14'd305,  -14'd467,  -14'd193,  -14'd1375,  -14'd1485,  14'd1426,  -14'd711,  
-14'd1552,  14'd1069,  14'd357,  -14'd1114,  14'd1490,  14'd145,  -14'd74,  14'd250,  14'd433,  -14'd288,  -14'd727,  14'd1411,  -14'd1059,  14'd498,  -14'd152,  -14'd998,  
14'd758,  14'd496,  14'd1997,  14'd569,  -14'd267,  14'd1641,  -14'd44,  14'd244,  14'd536,  14'd329,  14'd738,  14'd206,  14'd253,  14'd1069,  -14'd80,  -14'd404,  
14'd1081,  14'd115,  14'd132,  -14'd111,  -14'd1555,  14'd1406,  -14'd1204,  14'd1752,  14'd445,  14'd103,  -14'd673,  -14'd429,  14'd155,  14'd2619,  -14'd629,  -14'd213,  
-14'd101,  14'd108,  14'd388,  14'd1576,  14'd527,  14'd225,  -14'd1072,  14'd1163,  -14'd756,  14'd267,  -14'd304,  -14'd262,  14'd966,  14'd74,  14'd1001,  14'd30,  
14'd653,  -14'd705,  -14'd1029,  14'd724,  14'd470,  14'd1178,  14'd273,  14'd249,  -14'd632,  -14'd1361,  14'd1390,  14'd495,  14'd2002,  -14'd2312,  14'd235,  -14'd3,  
14'd1085,  14'd163,  -14'd228,  -14'd738,  -14'd185,  -14'd580,  14'd772,  14'd642,  14'd1283,  -14'd160,  14'd286,  14'd1356,  -14'd284,  -14'd270,  -14'd174,  -14'd1259,  
14'd1098,  -14'd685,  14'd456,  14'd193,  -14'd1236,  14'd428,  -14'd872,  -14'd1141,  14'd786,  -14'd181,  14'd275,  14'd1230,  14'd1462,  14'd1558,  -14'd1768,  14'd878,  

14'd194,  -14'd165,  -14'd1188,  14'd1059,  14'd603,  -14'd428,  -14'd292,  14'd75,  -14'd912,  14'd1349,  14'd660,  -14'd322,  -14'd97,  -14'd834,  14'd142,  14'd882,  
-14'd238,  -14'd1692,  -14'd310,  14'd721,  14'd471,  14'd675,  -14'd1074,  14'd1233,  14'd691,  -14'd118,  -14'd1530,  -14'd1114,  14'd1490,  -14'd913,  14'd375,  14'd62,  
-14'd1617,  -14'd279,  14'd939,  -14'd579,  14'd1102,  -14'd550,  -14'd45,  14'd721,  -14'd767,  14'd745,  14'd207,  14'd1070,  -14'd575,  -14'd882,  14'd86,  -14'd1299,  
-14'd1675,  -14'd2809,  14'd965,  -14'd1079,  -14'd344,  -14'd819,  14'd224,  -14'd642,  -14'd492,  -14'd534,  14'd1073,  14'd84,  -14'd1570,  14'd1410,  14'd1494,  -14'd1215,  
14'd163,  14'd415,  14'd288,  14'd554,  -14'd2009,  14'd445,  -14'd160,  14'd585,  14'd200,  -14'd535,  -14'd494,  14'd242,  -14'd1636,  14'd149,  14'd1434,  -14'd833,  
-14'd432,  14'd734,  -14'd177,  -14'd270,  -14'd111,  -14'd1040,  14'd16,  -14'd756,  14'd505,  -14'd2041,  14'd852,  14'd491,  14'd1173,  -14'd1414,  14'd720,  14'd996,  
-14'd454,  14'd2185,  14'd533,  14'd636,  14'd1312,  -14'd214,  14'd142,  -14'd849,  -14'd1259,  -14'd790,  -14'd685,  14'd407,  14'd123,  -14'd1639,  14'd697,  14'd1781,  
-14'd117,  -14'd635,  -14'd306,  14'd1095,  14'd678,  -14'd1078,  -14'd509,  14'd417,  14'd577,  14'd447,  -14'd1297,  14'd1261,  -14'd537,  14'd330,  14'd33,  14'd827,  
14'd440,  -14'd261,  14'd330,  14'd712,  -14'd140,  -14'd49,  -14'd173,  -14'd212,  14'd165,  -14'd329,  14'd1287,  14'd778,  14'd50,  -14'd1366,  14'd1142,  -14'd1853,  
14'd2179,  14'd847,  14'd968,  -14'd2,  14'd534,  14'd248,  14'd102,  -14'd987,  14'd368,  -14'd90,  -14'd545,  -14'd944,  14'd1481,  14'd844,  14'd571,  -14'd193,  
14'd179,  14'd843,  -14'd1,  -14'd897,  -14'd2385,  14'd770,  14'd668,  14'd56,  14'd1261,  14'd200,  14'd1470,  -14'd1059,  14'd651,  14'd335,  -14'd1162,  -14'd148,  
14'd250,  14'd1809,  -14'd122,  -14'd309,  14'd65,  14'd922,  -14'd235,  14'd1104,  14'd508,  14'd978,  -14'd1644,  14'd1803,  14'd354,  14'd459,  -14'd169,  -14'd288,  
-14'd599,  14'd1331,  14'd478,  -14'd474,  14'd427,  14'd473,  14'd27,  14'd1665,  -14'd494,  14'd747,  -14'd1043,  -14'd795,  14'd1433,  -14'd309,  14'd572,  -14'd1482,  
-14'd2833,  -14'd901,  -14'd445,  14'd160,  -14'd393,  14'd366,  -14'd1813,  -14'd65,  14'd120,  -14'd437,  -14'd1224,  14'd188,  14'd1181,  -14'd2495,  14'd782,  14'd1218,  
-14'd1041,  -14'd1559,  -14'd1218,  -14'd375,  14'd443,  -14'd1473,  14'd11,  14'd768,  14'd1120,  -14'd300,  -14'd506,  -14'd481,  14'd369,  14'd1198,  -14'd442,  -14'd52,  
14'd80,  -14'd902,  14'd1672,  14'd1452,  -14'd1146,  14'd1654,  14'd17,  14'd771,  14'd468,  14'd185,  14'd731,  -14'd971,  -14'd568,  14'd147,  14'd385,  -14'd1581,  
14'd1850,  14'd534,  -14'd829,  -14'd290,  -14'd593,  14'd71,  -14'd200,  14'd230,  -14'd581,  -14'd277,  -14'd275,  14'd625,  -14'd1344,  -14'd859,  14'd666,  -14'd581,  
14'd319,  14'd1731,  -14'd616,  -14'd393,  -14'd79,  14'd150,  -14'd522,  14'd601,  -14'd786,  -14'd751,  14'd917,  -14'd39,  -14'd856,  -14'd769,  14'd1462,  -14'd1593,  
-14'd416,  14'd532,  -14'd93,  14'd1190,  14'd1684,  14'd4,  -14'd831,  -14'd363,  14'd295,  -14'd718,  -14'd314,  14'd1604,  -14'd252,  14'd89,  14'd100,  -14'd313,  
-14'd571,  -14'd713,  14'd473,  14'd1457,  -14'd1036,  -14'd33,  -14'd9,  14'd3,  14'd505,  -14'd889,  -14'd52,  14'd272,  -14'd1245,  14'd1501,  14'd149,  14'd273,  
-14'd27,  -14'd194,  -14'd963,  -14'd873,  -14'd400,  14'd736,  14'd1104,  14'd224,  14'd639,  14'd1240,  14'd496,  -14'd39,  14'd345,  14'd315,  -14'd223,  -14'd862,  
14'd964,  14'd670,  -14'd1107,  -14'd1040,  14'd359,  -14'd267,  -14'd2110,  -14'd213,  14'd483,  14'd666,  14'd578,  14'd120,  -14'd1003,  -14'd1730,  14'd305,  -14'd599,  
14'd401,  -14'd420,  -14'd1125,  -14'd6,  14'd63,  14'd838,  -14'd460,  -14'd196,  -14'd32,  -14'd68,  14'd214,  14'd1648,  14'd502,  -14'd1445,  14'd899,  14'd38,  
14'd1714,  -14'd48,  14'd1758,  -14'd251,  -14'd837,  14'd160,  -14'd264,  14'd1107,  14'd2342,  14'd395,  14'd18,  14'd19,  -14'd803,  -14'd406,  -14'd491,  14'd179,  
14'd493,  14'd2633,  14'd1323,  14'd47,  -14'd1005,  -14'd1149,  14'd226,  -14'd465,  14'd1493,  -14'd2533,  -14'd245,  14'd314,  -14'd172,  14'd1057,  14'd210,  -14'd600,  

-14'd804,  -14'd389,  14'd169,  14'd88,  14'd431,  14'd407,  14'd831,  14'd338,  -14'd982,  14'd1433,  -14'd255,  14'd984,  14'd189,  14'd47,  14'd759,  -14'd907,  
14'd1043,  -14'd36,  -14'd1235,  14'd1442,  14'd2382,  14'd2282,  -14'd252,  14'd1387,  14'd983,  14'd1269,  -14'd50,  14'd681,  14'd474,  -14'd987,  -14'd368,  14'd93,  
14'd1286,  -14'd362,  -14'd103,  14'd220,  -14'd829,  -14'd335,  14'd1311,  14'd1148,  -14'd81,  -14'd354,  -14'd1137,  14'd648,  14'd909,  -14'd2235,  14'd798,  14'd782,  
14'd862,  14'd368,  -14'd176,  -14'd208,  14'd814,  14'd829,  14'd1550,  -14'd331,  -14'd1435,  -14'd1082,  14'd1198,  14'd987,  14'd2125,  14'd662,  14'd747,  14'd1138,  
-14'd594,  14'd613,  14'd142,  -14'd173,  14'd685,  -14'd505,  14'd1156,  -14'd310,  14'd297,  14'd1087,  -14'd542,  14'd246,  -14'd1044,  14'd469,  14'd1104,  -14'd995,  
-14'd116,  14'd1233,  14'd477,  14'd1491,  -14'd408,  -14'd1132,  -14'd721,  -14'd611,  -14'd861,  -14'd883,  14'd2251,  14'd172,  14'd173,  14'd1514,  14'd690,  14'd248,  
14'd700,  14'd1664,  -14'd364,  14'd611,  14'd2245,  -14'd757,  14'd268,  -14'd1451,  14'd596,  -14'd511,  14'd469,  14'd746,  -14'd513,  -14'd2649,  -14'd1213,  14'd705,  
14'd290,  14'd331,  -14'd400,  -14'd1283,  14'd244,  -14'd1229,  14'd927,  -14'd798,  14'd2423,  14'd826,  14'd887,  14'd1302,  -14'd753,  -14'd535,  -14'd755,  14'd2313,  
14'd1333,  14'd843,  14'd197,  14'd312,  -14'd584,  -14'd786,  14'd194,  -14'd861,  14'd956,  -14'd269,  14'd1835,  -14'd812,  14'd943,  -14'd782,  14'd186,  -14'd44,  
-14'd679,  14'd1424,  -14'd1588,  14'd29,  -14'd1417,  14'd882,  14'd56,  -14'd639,  14'd1438,  -14'd1559,  14'd853,  -14'd2062,  14'd97,  14'd1805,  14'd297,  14'd514,  
14'd314,  14'd669,  14'd1356,  14'd535,  -14'd2908,  14'd250,  14'd1504,  14'd226,  14'd114,  -14'd686,  14'd949,  -14'd1237,  -14'd64,  -14'd329,  -14'd413,  14'd1150,  
14'd435,  14'd1068,  -14'd1333,  -14'd2149,  -14'd117,  14'd251,  -14'd307,  -14'd1257,  -14'd510,  -14'd840,  -14'd743,  -14'd256,  -14'd1953,  14'd1094,  -14'd1113,  14'd398,  
14'd525,  14'd1308,  -14'd202,  -14'd1172,  -14'd531,  -14'd541,  -14'd304,  14'd437,  -14'd760,  14'd1196,  -14'd602,  -14'd1528,  14'd505,  14'd2214,  14'd998,  -14'd1207,  
-14'd12,  14'd393,  -14'd562,  -14'd335,  14'd1658,  -14'd358,  -14'd500,  -14'd381,  -14'd758,  14'd480,  -14'd6,  -14'd153,  -14'd760,  14'd492,  14'd657,  -14'd747,  
-14'd1684,  14'd409,  14'd13,  -14'd497,  14'd1332,  14'd411,  -14'd430,  14'd614,  -14'd509,  14'd137,  -14'd1227,  -14'd1097,  -14'd1088,  14'd1644,  14'd1574,  14'd1061,  
14'd179,  -14'd2045,  14'd58,  -14'd1801,  -14'd661,  -14'd26,  14'd439,  -14'd265,  14'd875,  14'd832,  -14'd74,  -14'd1201,  -14'd84,  14'd517,  -14'd2056,  -14'd1667,  
14'd447,  14'd1251,  14'd1194,  -14'd181,  -14'd1729,  -14'd583,  14'd1102,  -14'd423,  -14'd1330,  14'd130,  -14'd587,  -14'd875,  -14'd420,  14'd578,  14'd434,  -14'd1159,  
-14'd852,  -14'd886,  14'd519,  -14'd1840,  14'd484,  14'd605,  14'd1120,  14'd263,  14'd287,  -14'd413,  14'd585,  14'd359,  -14'd1293,  14'd486,  -14'd823,  14'd1079,  
-14'd2458,  -14'd715,  -14'd2359,  14'd993,  14'd1513,  14'd1070,  14'd83,  -14'd966,  14'd263,  -14'd1829,  -14'd1263,  -14'd230,  -14'd924,  -14'd499,  14'd953,  -14'd404,  
-14'd543,  14'd537,  14'd954,  -14'd220,  14'd415,  14'd1000,  14'd809,  -14'd1487,  14'd918,  -14'd733,  -14'd870,  14'd736,  -14'd1330,  -14'd487,  14'd1070,  -14'd475,  
-14'd1432,  -14'd216,  14'd428,  14'd1516,  14'd764,  14'd317,  14'd1639,  14'd951,  14'd1373,  14'd556,  -14'd1252,  -14'd443,  14'd834,  14'd501,  14'd1435,  -14'd768,  
14'd659,  14'd198,  14'd361,  14'd199,  -14'd408,  -14'd625,  -14'd1433,  14'd170,  -14'd403,  14'd1086,  -14'd976,  14'd813,  -14'd1523,  -14'd1780,  14'd66,  -14'd581,  
-14'd105,  -14'd412,  -14'd2,  -14'd1085,  -14'd370,  14'd361,  -14'd854,  -14'd105,  -14'd509,  14'd1783,  -14'd851,  14'd674,  -14'd950,  -14'd824,  -14'd533,  14'd533,  
14'd743,  14'd1089,  14'd1093,  -14'd846,  -14'd635,  14'd511,  -14'd383,  -14'd424,  14'd362,  14'd691,  -14'd1438,  14'd158,  -14'd85,  14'd617,  -14'd313,  -14'd916,  
14'd2672,  14'd1071,  14'd3111,  14'd1898,  -14'd1770,  14'd2058,  14'd55,  -14'd65,  14'd1967,  -14'd1206,  -14'd678,  14'd642,  14'd1192,  -14'd83,  -14'd1064,  -14'd958,  

14'd76,  -14'd931,  -14'd1251,  14'd27,  -14'd691,  14'd225,  -14'd307,  -14'd126,  14'd885,  -14'd839,  14'd546,  -14'd108,  -14'd407,  -14'd300,  -14'd249,  -14'd445,  
-14'd1288,  14'd1097,  14'd124,  -14'd1949,  14'd183,  -14'd1222,  14'd527,  -14'd769,  14'd733,  14'd24,  14'd65,  -14'd1017,  14'd243,  -14'd35,  -14'd816,  14'd403,  
14'd553,  14'd52,  -14'd159,  -14'd799,  14'd455,  -14'd1131,  -14'd917,  -14'd138,  -14'd386,  -14'd155,  -14'd382,  -14'd903,  -14'd1444,  -14'd219,  -14'd122,  -14'd1017,  
14'd798,  -14'd863,  -14'd502,  -14'd1022,  -14'd155,  -14'd472,  14'd246,  -14'd582,  -14'd1155,  -14'd266,  -14'd1484,  14'd264,  -14'd665,  -14'd1514,  -14'd196,  14'd147,  
-14'd29,  -14'd1042,  14'd62,  14'd1146,  -14'd216,  14'd1158,  -14'd1696,  14'd1135,  -14'd757,  14'd730,  14'd363,  -14'd236,  -14'd1006,  14'd406,  -14'd105,  14'd250,  
14'd674,  -14'd886,  14'd716,  14'd890,  -14'd1381,  14'd187,  14'd785,  -14'd822,  -14'd1530,  -14'd879,  14'd444,  -14'd606,  -14'd524,  14'd542,  14'd82,  14'd509,  
-14'd235,  -14'd870,  -14'd154,  -14'd104,  -14'd1379,  -14'd277,  -14'd343,  -14'd107,  -14'd249,  -14'd950,  -14'd490,  -14'd1015,  14'd352,  14'd852,  14'd373,  -14'd700,  
-14'd1551,  -14'd49,  -14'd733,  -14'd684,  -14'd801,  -14'd241,  -14'd602,  -14'd908,  -14'd1046,  -14'd1017,  -14'd591,  14'd758,  14'd276,  -14'd310,  -14'd1684,  14'd595,  
-14'd653,  -14'd221,  -14'd374,  14'd198,  14'd794,  -14'd670,  -14'd292,  -14'd465,  -14'd1058,  -14'd554,  14'd403,  14'd848,  -14'd188,  -14'd316,  14'd170,  -14'd482,  
14'd121,  -14'd864,  -14'd756,  -14'd918,  -14'd482,  -14'd284,  -14'd764,  14'd324,  14'd317,  -14'd678,  -14'd900,  14'd258,  14'd990,  14'd825,  14'd631,  -14'd457,  
-14'd1494,  14'd146,  -14'd28,  -14'd764,  14'd353,  14'd188,  -14'd531,  -14'd307,  14'd281,  -14'd230,  -14'd857,  14'd180,  14'd328,  14'd379,  -14'd509,  -14'd1381,  
-14'd351,  -14'd1232,  14'd35,  -14'd1649,  -14'd1156,  14'd337,  14'd690,  -14'd460,  -14'd425,  14'd310,  14'd1088,  -14'd36,  14'd541,  14'd318,  -14'd1811,  -14'd1562,  
14'd323,  -14'd1546,  14'd1281,  -14'd36,  -14'd1092,  -14'd1279,  14'd389,  -14'd103,  -14'd1047,  14'd805,  -14'd479,  14'd580,  14'd38,  14'd1187,  14'd60,  -14'd1117,  
14'd1398,  14'd172,  14'd45,  -14'd1368,  -14'd855,  -14'd379,  -14'd293,  -14'd714,  -14'd90,  14'd603,  14'd662,  -14'd502,  -14'd212,  -14'd799,  14'd508,  14'd208,  
-14'd313,  -14'd10,  14'd248,  14'd817,  -14'd468,  -14'd842,  -14'd1164,  -14'd663,  -14'd372,  -14'd69,  -14'd284,  14'd1058,  14'd312,  -14'd369,  14'd477,  -14'd233,  
14'd1300,  -14'd1549,  -14'd922,  14'd384,  -14'd1779,  14'd185,  14'd613,  -14'd1183,  -14'd267,  -14'd952,  14'd723,  14'd313,  -14'd464,  -14'd764,  -14'd794,  -14'd245,  
14'd233,  14'd463,  14'd369,  14'd732,  -14'd418,  -14'd1352,  14'd890,  14'd636,  -14'd418,  14'd240,  -14'd574,  14'd471,  14'd221,  -14'd1116,  -14'd169,  -14'd787,  
-14'd577,  -14'd416,  -14'd307,  -14'd1173,  -14'd339,  -14'd431,  14'd419,  -14'd268,  -14'd115,  -14'd250,  14'd1045,  -14'd1109,  -14'd218,  -14'd36,  -14'd846,  14'd467,  
-14'd1151,  14'd859,  14'd1101,  14'd80,  14'd391,  -14'd720,  -14'd1359,  -14'd543,  -14'd956,  -14'd1299,  14'd583,  -14'd747,  14'd62,  14'd188,  14'd984,  14'd300,  
-14'd834,  -14'd879,  -14'd1003,  -14'd1225,  -14'd635,  14'd619,  14'd881,  14'd6,  -14'd1310,  14'd321,  14'd587,  14'd1127,  -14'd470,  -14'd1093,  14'd140,  -14'd249,  
14'd407,  -14'd1089,  14'd437,  -14'd695,  -14'd804,  -14'd971,  14'd555,  14'd534,  -14'd254,  -14'd767,  -14'd146,  14'd853,  -14'd99,  -14'd396,  14'd306,  -14'd148,  
-14'd509,  -14'd1739,  -14'd71,  14'd25,  -14'd237,  14'd565,  -14'd923,  -14'd1553,  -14'd226,  -14'd282,  14'd628,  -14'd701,  14'd112,  14'd82,  -14'd1456,  -14'd119,  
-14'd702,  -14'd460,  14'd1013,  14'd391,  14'd976,  -14'd378,  -14'd1073,  -14'd328,  14'd68,  -14'd447,  14'd1198,  -14'd1348,  -14'd1240,  -14'd18,  14'd264,  -14'd1380,  
-14'd466,  -14'd40,  14'd690,  -14'd174,  14'd751,  14'd391,  -14'd648,  14'd178,  -14'd180,  14'd11,  14'd398,  -14'd189,  -14'd1075,  -14'd1648,  -14'd29,  14'd198,  
-14'd1115,  -14'd17,  -14'd331,  -14'd601,  14'd101,  -14'd1387,  14'd840,  14'd404,  -14'd1288,  14'd65,  -14'd8,  -14'd2047,  14'd275,  14'd342,  -14'd501,  14'd199,  

14'd344,  -14'd833,  14'd656,  -14'd1684,  -14'd496,  -14'd714,  14'd1460,  -14'd58,  14'd66,  -14'd186,  -14'd1577,  -14'd201,  -14'd479,  14'd348,  -14'd242,  -14'd273,  
14'd1772,  14'd1167,  -14'd104,  -14'd1517,  -14'd1708,  14'd1855,  14'd2142,  14'd387,  14'd267,  -14'd106,  -14'd185,  -14'd1,  14'd1360,  14'd2091,  14'd94,  -14'd113,  
14'd283,  -14'd562,  -14'd425,  14'd317,  -14'd308,  14'd519,  14'd1653,  -14'd55,  14'd258,  -14'd823,  14'd1140,  14'd439,  14'd235,  14'd740,  14'd4,  14'd742,  
14'd951,  14'd984,  14'd434,  14'd273,  14'd1951,  14'd2375,  -14'd873,  14'd444,  14'd1982,  14'd276,  14'd218,  -14'd620,  14'd791,  -14'd368,  14'd979,  -14'd32,  
14'd686,  14'd197,  14'd94,  -14'd1234,  14'd51,  -14'd190,  -14'd386,  14'd1387,  -14'd1427,  14'd134,  14'd1265,  14'd393,  14'd1875,  -14'd805,  14'd399,  -14'd349,  
-14'd184,  -14'd1821,  14'd595,  -14'd1124,  -14'd20,  14'd674,  14'd1008,  -14'd44,  -14'd756,  -14'd13,  14'd966,  -14'd542,  -14'd1433,  14'd0,  14'd160,  14'd93,  
-14'd211,  14'd212,  14'd1000,  -14'd1434,  14'd1207,  14'd110,  14'd789,  14'd501,  -14'd313,  -14'd117,  14'd1842,  14'd565,  14'd879,  14'd858,  -14'd496,  -14'd220,  
14'd457,  -14'd180,  14'd1891,  -14'd93,  -14'd452,  14'd1248,  14'd472,  14'd730,  14'd627,  -14'd331,  -14'd30,  -14'd1703,  -14'd473,  -14'd184,  14'd459,  -14'd979,  
14'd1052,  14'd1099,  -14'd39,  -14'd756,  -14'd40,  14'd961,  -14'd1869,  -14'd516,  14'd246,  -14'd247,  14'd582,  -14'd93,  14'd378,  -14'd1003,  -14'd1490,  14'd1128,  
-14'd1731,  -14'd968,  14'd2233,  14'd627,  -14'd817,  14'd159,  -14'd92,  -14'd734,  -14'd37,  14'd563,  14'd5,  14'd1546,  -14'd306,  -14'd490,  14'd1191,  14'd1838,  
-14'd913,  14'd1519,  -14'd282,  -14'd475,  -14'd1832,  -14'd1697,  14'd555,  14'd40,  -14'd2735,  -14'd862,  -14'd1210,  14'd5,  -14'd1040,  14'd335,  14'd1088,  14'd420,  
14'd1312,  -14'd1310,  14'd176,  -14'd475,  -14'd1008,  -14'd1292,  -14'd817,  -14'd1788,  -14'd756,  -14'd1638,  -14'd5,  14'd799,  -14'd1456,  14'd716,  -14'd6,  14'd92,  
-14'd313,  -14'd159,  -14'd40,  14'd105,  -14'd455,  -14'd848,  -14'd5,  14'd246,  14'd687,  -14'd968,  -14'd372,  -14'd445,  -14'd1195,  -14'd833,  14'd709,  14'd15,  
-14'd2100,  14'd787,  -14'd657,  -14'd717,  14'd1326,  -14'd747,  14'd1134,  -14'd931,  -14'd588,  14'd650,  14'd131,  14'd392,  -14'd681,  -14'd394,  -14'd614,  -14'd781,  
-14'd971,  -14'd322,  14'd914,  -14'd302,  -14'd1186,  14'd1677,  14'd317,  -14'd82,  -14'd364,  14'd193,  -14'd126,  14'd535,  -14'd3632,  -14'd170,  -14'd408,  14'd62,  
14'd595,  14'd748,  14'd1450,  -14'd1054,  -14'd1175,  -14'd408,  14'd702,  14'd348,  -14'd2100,  -14'd939,  -14'd1746,  14'd86,  14'd7,  14'd1291,  -14'd158,  14'd875,  
14'd1044,  -14'd17,  14'd2223,  -14'd772,  -14'd407,  14'd1347,  14'd1935,  14'd1178,  14'd223,  -14'd1585,  -14'd1008,  14'd412,  -14'd1676,  14'd2028,  14'd977,  14'd130,  
14'd229,  -14'd53,  -14'd1383,  14'd49,  -14'd108,  -14'd1230,  14'd688,  14'd456,  -14'd1623,  -14'd761,  -14'd316,  14'd211,  -14'd2349,  14'd329,  -14'd750,  -14'd871,  
-14'd1597,  -14'd257,  -14'd1019,  14'd472,  -14'd598,  -14'd448,  -14'd254,  -14'd722,  -14'd553,  -14'd431,  -14'd1282,  14'd595,  14'd807,  14'd1403,  14'd326,  -14'd676,  
-14'd203,  -14'd163,  -14'd329,  -14'd1248,  14'd404,  14'd541,  14'd1040,  -14'd631,  14'd2225,  14'd534,  -14'd522,  -14'd987,  -14'd1622,  14'd557,  -14'd662,  -14'd2150,  
-14'd125,  -14'd1050,  14'd529,  -14'd531,  -14'd264,  14'd54,  14'd184,  14'd459,  -14'd1723,  14'd1374,  -14'd1166,  -14'd1175,  -14'd246,  14'd2025,  -14'd272,  -14'd225,  
-14'd1,  -14'd813,  14'd379,  14'd1660,  14'd877,  14'd1889,  -14'd1034,  14'd220,  -14'd456,  -14'd31,  -14'd186,  -14'd310,  -14'd572,  -14'd1044,  14'd1556,  14'd306,  
-14'd520,  14'd842,  -14'd1106,  14'd1171,  -14'd480,  -14'd173,  14'd411,  -14'd256,  14'd572,  14'd324,  -14'd177,  -14'd1127,  14'd512,  14'd236,  14'd812,  -14'd1504,  
-14'd1076,  -14'd703,  -14'd29,  -14'd744,  14'd1533,  -14'd1773,  14'd265,  -14'd149,  14'd1382,  14'd42,  14'd518,  14'd819,  -14'd17,  14'd121,  14'd113,  -14'd189,  
14'd731,  -14'd760,  -14'd940,  14'd1122,  -14'd55,  14'd1431,  -14'd574,  -14'd796,  14'd969,  14'd1757,  -14'd1497,  14'd1551,  14'd619,  -14'd49,  14'd9,  -14'd442,  

-14'd2055,  14'd22,  -14'd696,  -14'd38,  14'd1638,  14'd441,  -14'd521,  -14'd179,  14'd235,  -14'd1027,  14'd261,  14'd659,  14'd1357,  -14'd542,  14'd121,  14'd999,  
14'd14,  14'd739,  -14'd93,  -14'd52,  14'd2027,  -14'd742,  14'd434,  14'd37,  14'd1219,  -14'd986,  -14'd905,  14'd1065,  -14'd84,  14'd726,  -14'd30,  14'd394,  
-14'd168,  14'd1650,  14'd127,  -14'd1787,  14'd58,  -14'd7,  14'd377,  -14'd164,  -14'd1357,  -14'd1050,  -14'd1203,  -14'd56,  -14'd745,  14'd2711,  -14'd16,  14'd933,  
-14'd1020,  14'd1223,  -14'd406,  14'd391,  14'd260,  14'd507,  14'd1739,  -14'd49,  14'd411,  14'd318,  14'd123,  -14'd1299,  -14'd598,  14'd3185,  14'd132,  14'd745,  
-14'd236,  14'd607,  -14'd508,  -14'd1423,  14'd417,  14'd469,  14'd984,  14'd1037,  14'd1185,  14'd1356,  14'd850,  -14'd604,  -14'd1403,  14'd1212,  14'd847,  -14'd1192,  
-14'd656,  14'd237,  14'd496,  14'd24,  14'd366,  -14'd876,  14'd2440,  -14'd690,  -14'd587,  -14'd711,  14'd973,  14'd863,  14'd827,  -14'd327,  -14'd1464,  14'd902,  
14'd298,  14'd144,  -14'd448,  -14'd127,  14'd263,  -14'd25,  14'd311,  -14'd106,  -14'd329,  14'd1105,  -14'd246,  14'd685,  -14'd698,  -14'd206,  -14'd440,  -14'd445,  
14'd267,  -14'd984,  -14'd156,  -14'd1604,  -14'd485,  -14'd778,  14'd244,  -14'd488,  -14'd437,  14'd961,  -14'd1391,  14'd773,  -14'd755,  -14'd745,  -14'd592,  -14'd1601,  
-14'd665,  -14'd1379,  14'd1820,  14'd857,  -14'd306,  14'd695,  14'd829,  -14'd1825,  -14'd859,  14'd598,  14'd1425,  14'd221,  14'd356,  14'd1,  -14'd228,  -14'd801,  
14'd863,  14'd1454,  14'd646,  14'd354,  -14'd1345,  14'd386,  14'd101,  -14'd529,  14'd724,  14'd513,  -14'd20,  14'd416,  14'd487,  -14'd1512,  14'd109,  -14'd252,  
14'd951,  14'd870,  14'd217,  -14'd1501,  -14'd1553,  14'd168,  14'd511,  -14'd797,  -14'd662,  14'd681,  14'd1818,  14'd857,  -14'd1104,  -14'd546,  -14'd996,  14'd3,  
-14'd363,  14'd927,  -14'd935,  14'd1326,  14'd518,  14'd1634,  -14'd250,  14'd217,  14'd970,  -14'd1072,  -14'd441,  14'd1035,  14'd243,  -14'd189,  14'd1031,  14'd1517,  
-14'd107,  14'd660,  14'd667,  -14'd266,  -14'd505,  14'd310,  14'd40,  -14'd205,  14'd767,  14'd1200,  14'd130,  -14'd247,  14'd737,  14'd883,  -14'd193,  14'd221,  
-14'd627,  14'd29,  14'd914,  14'd795,  -14'd992,  -14'd401,  -14'd446,  -14'd1704,  14'd69,  14'd625,  14'd247,  14'd119,  14'd460,  14'd447,  -14'd290,  14'd1455,  
14'd1229,  -14'd842,  14'd241,  14'd1284,  -14'd310,  14'd931,  14'd824,  -14'd403,  14'd425,  14'd659,  14'd1087,  14'd740,  14'd331,  -14'd715,  -14'd1438,  -14'd1006,  
14'd1233,  14'd925,  -14'd178,  -14'd588,  -14'd2074,  14'd700,  14'd744,  -14'd376,  -14'd1428,  -14'd1504,  14'd144,  14'd2070,  14'd1117,  14'd582,  14'd649,  14'd1625,  
14'd2298,  -14'd1301,  14'd298,  14'd159,  14'd499,  14'd363,  14'd152,  -14'd148,  14'd841,  14'd680,  14'd203,  14'd327,  -14'd875,  14'd490,  14'd1648,  -14'd921,  
14'd528,  14'd186,  -14'd1175,  14'd1047,  14'd674,  -14'd279,  -14'd406,  14'd661,  14'd451,  14'd365,  14'd26,  14'd999,  14'd1578,  -14'd1064,  -14'd845,  14'd1193,  
14'd435,  14'd484,  -14'd266,  -14'd446,  14'd1190,  -14'd1336,  -14'd1753,  -14'd733,  14'd235,  14'd76,  14'd312,  -14'd1219,  14'd559,  -14'd870,  14'd437,  14'd441,  
14'd920,  14'd1000,  14'd532,  -14'd368,  14'd436,  14'd84,  -14'd404,  14'd484,  14'd529,  -14'd302,  14'd1356,  14'd778,  14'd13,  14'd599,  -14'd821,  14'd1344,  
14'd1676,  14'd1,  14'd457,  14'd1797,  14'd784,  14'd353,  -14'd59,  14'd956,  -14'd700,  14'd1681,  -14'd237,  14'd434,  14'd814,  14'd1377,  14'd64,  14'd916,  
14'd386,  -14'd386,  14'd589,  -14'd172,  14'd851,  14'd960,  -14'd1155,  14'd1518,  -14'd2534,  -14'd495,  14'd1208,  -14'd896,  14'd389,  14'd966,  -14'd930,  14'd45,  
14'd560,  -14'd236,  -14'd482,  14'd509,  -14'd963,  14'd1456,  14'd739,  14'd1278,  -14'd2137,  -14'd312,  -14'd279,  -14'd338,  14'd359,  -14'd1933,  14'd562,  14'd754,  
14'd364,  -14'd143,  -14'd579,  -14'd305,  14'd1215,  -14'd1282,  -14'd324,  14'd546,  -14'd434,  14'd120,  -14'd445,  -14'd1205,  14'd1334,  -14'd19,  14'd737,  -14'd775,  
14'd302,  -14'd876,  -14'd1964,  -14'd73,  14'd991,  14'd824,  14'd623,  14'd648,  -14'd937,  -14'd307,  14'd501,  14'd1298,  14'd1668,  -14'd733,  -14'd881,  14'd296,  

14'd2116,  14'd557,  14'd1311,  14'd1520,  -14'd453,  14'd949,  14'd2311,  14'd1557,  -14'd90,  -14'd923,  14'd361,  -14'd571,  14'd318,  14'd2160,  -14'd200,  -14'd801,  
-14'd25,  14'd693,  14'd465,  14'd1638,  -14'd1056,  14'd759,  -14'd283,  -14'd133,  14'd749,  -14'd418,  14'd1065,  14'd2095,  14'd112,  14'd889,  14'd86,  14'd1046,  
-14'd765,  14'd280,  14'd443,  14'd586,  14'd1144,  -14'd460,  14'd1031,  -14'd108,  14'd1416,  14'd2165,  14'd1609,  14'd247,  14'd562,  14'd972,  -14'd937,  -14'd298,  
-14'd1088,  -14'd800,  14'd2628,  14'd68,  -14'd810,  -14'd315,  -14'd1438,  14'd1367,  -14'd209,  14'd1304,  -14'd639,  14'd1054,  14'd527,  14'd1409,  14'd1234,  14'd136,  
-14'd856,  -14'd2770,  -14'd812,  -14'd648,  -14'd183,  -14'd1318,  -14'd1257,  -14'd782,  -14'd2600,  14'd401,  14'd457,  -14'd302,  -14'd6,  -14'd372,  -14'd910,  -14'd956,  
14'd504,  -14'd357,  14'd1444,  14'd970,  -14'd1558,  -14'd107,  -14'd807,  -14'd291,  14'd316,  14'd1134,  -14'd295,  14'd268,  14'd993,  14'd132,  14'd229,  14'd706,  
-14'd546,  -14'd186,  14'd1606,  14'd1643,  -14'd1131,  14'd702,  14'd602,  14'd917,  -14'd977,  14'd1042,  14'd607,  -14'd1410,  14'd1167,  -14'd574,  14'd119,  14'd420,  
-14'd29,  14'd116,  -14'd1368,  14'd1221,  -14'd146,  14'd240,  -14'd1262,  14'd389,  -14'd1274,  -14'd1117,  -14'd386,  -14'd579,  14'd1792,  14'd434,  14'd1204,  14'd613,  
-14'd988,  14'd660,  14'd716,  14'd943,  -14'd2050,  14'd318,  -14'd865,  14'd257,  -14'd1381,  -14'd423,  -14'd994,  14'd79,  -14'd1956,  14'd1661,  14'd284,  -14'd728,  
-14'd366,  -14'd1767,  14'd1142,  -14'd158,  -14'd1958,  -14'd58,  -14'd1628,  14'd783,  -14'd623,  14'd556,  14'd726,  14'd724,  -14'd2033,  14'd1420,  -14'd343,  -14'd1969,  
14'd701,  14'd89,  -14'd1286,  -14'd867,  14'd322,  14'd133,  14'd1023,  -14'd151,  -14'd1210,  -14'd196,  14'd2383,  -14'd1308,  14'd741,  14'd331,  14'd302,  -14'd957,  
-14'd935,  14'd648,  -14'd1237,  -14'd381,  -14'd1314,  -14'd656,  -14'd2403,  -14'd274,  14'd250,  14'd299,  -14'd727,  -14'd1661,  14'd606,  -14'd183,  14'd920,  -14'd471,  
-14'd1204,  14'd1032,  -14'd1184,  14'd338,  14'd694,  -14'd1518,  14'd532,  -14'd1226,  14'd463,  -14'd1014,  -14'd793,  -14'd487,  -14'd678,  14'd913,  -14'd440,  -14'd417,  
-14'd1684,  14'd553,  14'd980,  -14'd554,  -14'd2113,  -14'd880,  -14'd442,  -14'd173,  -14'd1392,  -14'd887,  14'd2405,  14'd581,  -14'd1376,  -14'd470,  -14'd582,  -14'd701,  
14'd1050,  14'd507,  14'd331,  -14'd154,  14'd417,  -14'd96,  -14'd697,  -14'd1380,  -14'd1123,  -14'd1840,  -14'd229,  -14'd222,  -14'd786,  -14'd995,  14'd83,  -14'd335,  
-14'd139,  14'd133,  -14'd37,  -14'd1272,  -14'd879,  -14'd1353,  14'd724,  -14'd459,  14'd194,  -14'd179,  14'd48,  14'd99,  14'd450,  -14'd374,  -14'd232,  -14'd270,  
-14'd1432,  -14'd634,  14'd1204,  14'd270,  -14'd48,  -14'd1059,  -14'd204,  -14'd935,  14'd518,  14'd571,  14'd624,  14'd2121,  -14'd841,  -14'd756,  14'd894,  14'd1014,  
14'd116,  14'd217,  14'd1454,  14'd341,  14'd827,  14'd1396,  14'd1262,  -14'd71,  14'd2540,  14'd2447,  -14'd1908,  -14'd166,  -14'd399,  14'd1472,  14'd599,  -14'd2040,  
14'd439,  14'd87,  14'd1284,  14'd355,  -14'd598,  14'd346,  14'd292,  14'd32,  14'd434,  14'd220,  -14'd1182,  14'd532,  -14'd1061,  14'd629,  14'd949,  -14'd2177,  
14'd1444,  -14'd1127,  -14'd95,  -14'd126,  -14'd269,  -14'd413,  -14'd1156,  -14'd681,  14'd657,  14'd1021,  -14'd844,  14'd84,  14'd1189,  -14'd358,  14'd737,  -14'd543,  
14'd820,  -14'd303,  14'd113,  14'd1403,  -14'd800,  14'd173,  14'd1764,  14'd898,  -14'd86,  -14'd1308,  -14'd122,  14'd21,  -14'd70,  -14'd781,  -14'd16,  -14'd166,  
-14'd1015,  -14'd240,  14'd508,  14'd2050,  -14'd812,  14'd2115,  14'd269,  -14'd275,  14'd1751,  -14'd126,  14'd284,  14'd1042,  14'd702,  14'd636,  -14'd881,  14'd207,  
14'd674,  -14'd273,  14'd170,  14'd1777,  14'd1950,  14'd1355,  14'd610,  -14'd326,  -14'd881,  14'd428,  14'd1254,  -14'd848,  14'd1265,  14'd498,  -14'd55,  14'd325,  
-14'd1303,  14'd995,  -14'd1924,  14'd1334,  14'd360,  14'd267,  -14'd1029,  -14'd40,  14'd528,  14'd916,  14'd545,  -14'd611,  14'd915,  -14'd1483,  14'd1020,  14'd199,  
-14'd1482,  -14'd1356,  14'd281,  14'd1242,  14'd257,  14'd19,  -14'd427,  -14'd494,  -14'd425,  14'd2219,  14'd1359,  14'd507,  14'd853,  -14'd2255,  14'd860,  -14'd308,  

-14'd988,  14'd132,  14'd802,  14'd1305,  -14'd933,  -14'd190,  -14'd952,  14'd589,  -14'd558,  14'd569,  -14'd526,  -14'd1755,  14'd1896,  -14'd631,  14'd1255,  14'd214,  
14'd67,  -14'd291,  14'd208,  14'd175,  14'd329,  -14'd1286,  -14'd1078,  -14'd0,  14'd973,  -14'd26,  14'd48,  14'd1276,  -14'd565,  -14'd242,  14'd528,  -14'd90,  
14'd171,  -14'd280,  14'd1156,  14'd336,  14'd287,  -14'd614,  -14'd182,  14'd292,  -14'd371,  14'd220,  14'd281,  14'd196,  14'd1292,  14'd1324,  -14'd407,  -14'd1323,  
-14'd35,  14'd52,  -14'd756,  -14'd798,  14'd90,  -14'd589,  14'd66,  -14'd672,  -14'd65,  -14'd697,  -14'd602,  14'd215,  -14'd587,  14'd150,  -14'd428,  -14'd1125,  
14'd1286,  14'd734,  -14'd385,  14'd90,  -14'd610,  14'd116,  -14'd515,  -14'd539,  -14'd1110,  -14'd546,  14'd225,  14'd1372,  -14'd956,  14'd97,  -14'd211,  -14'd386,  
-14'd73,  14'd720,  14'd4,  14'd438,  14'd710,  14'd1300,  -14'd1283,  -14'd611,  14'd267,  14'd291,  -14'd233,  14'd1372,  -14'd385,  -14'd584,  14'd730,  -14'd649,  
-14'd413,  -14'd327,  14'd583,  14'd470,  14'd1340,  -14'd799,  14'd72,  14'd369,  14'd573,  -14'd646,  -14'd679,  14'd809,  14'd1181,  -14'd502,  14'd249,  -14'd309,  
-14'd776,  14'd484,  -14'd808,  14'd1275,  -14'd153,  -14'd395,  14'd684,  -14'd1575,  14'd387,  -14'd309,  14'd404,  -14'd1,  14'd996,  14'd1311,  -14'd238,  14'd578,  
-14'd387,  -14'd420,  -14'd113,  -14'd179,  14'd1812,  14'd139,  14'd286,  -14'd123,  14'd1877,  -14'd452,  14'd303,  -14'd341,  14'd51,  -14'd311,  -14'd171,  -14'd1259,  
14'd2845,  14'd327,  -14'd1209,  14'd1507,  14'd1319,  14'd530,  -14'd187,  14'd243,  -14'd66,  14'd1353,  -14'd156,  14'd268,  14'd1866,  14'd622,  14'd250,  14'd88,  
-14'd1134,  14'd488,  -14'd272,  14'd565,  14'd520,  14'd1380,  -14'd643,  14'd612,  14'd97,  -14'd971,  14'd93,  -14'd795,  -14'd294,  14'd134,  14'd996,  14'd961,  
-14'd279,  -14'd148,  -14'd48,  14'd406,  14'd212,  -14'd514,  -14'd495,  14'd1656,  -14'd1325,  14'd644,  -14'd920,  14'd1394,  14'd1059,  -14'd1668,  14'd720,  14'd1205,  
-14'd1312,  14'd611,  -14'd771,  14'd759,  -14'd858,  14'd743,  14'd1569,  -14'd484,  14'd365,  -14'd480,  14'd1668,  -14'd322,  14'd2175,  14'd119,  -14'd906,  -14'd189,  
-14'd432,  -14'd1018,  -14'd702,  14'd1646,  -14'd385,  14'd1040,  -14'd171,  -14'd224,  14'd1210,  -14'd20,  14'd1451,  -14'd1,  14'd1311,  -14'd601,  -14'd297,  14'd650,  
-14'd1870,  -14'd276,  14'd17,  14'd356,  -14'd169,  14'd558,  -14'd1614,  14'd713,  14'd567,  -14'd700,  14'd344,  -14'd1011,  14'd1215,  14'd385,  14'd916,  -14'd604,  
-14'd661,  14'd1099,  -14'd671,  -14'd892,  14'd1309,  -14'd1240,  -14'd1780,  -14'd747,  -14'd194,  14'd2038,  14'd1238,  -14'd1089,  -14'd800,  14'd618,  -14'd1782,  -14'd586,  
14'd203,  14'd1660,  -14'd654,  -14'd448,  -14'd339,  14'd643,  -14'd707,  14'd488,  14'd221,  14'd823,  14'd971,  -14'd1260,  14'd756,  -14'd3192,  -14'd1262,  -14'd405,  
-14'd258,  14'd779,  -14'd1717,  -14'd1331,  14'd786,  -14'd356,  14'd177,  -14'd897,  14'd656,  -14'd203,  14'd322,  -14'd1407,  -14'd418,  -14'd1139,  -14'd760,  14'd1510,  
-14'd1339,  14'd1323,  -14'd270,  -14'd854,  14'd1848,  -14'd656,  14'd1500,  -14'd931,  14'd1874,  14'd581,  -14'd18,  14'd1063,  -14'd170,  -14'd669,  14'd1050,  14'd1249,  
-14'd1030,  14'd458,  -14'd1970,  14'd266,  14'd57,  -14'd141,  14'd714,  14'd1156,  -14'd301,  -14'd1061,  14'd23,  14'd314,  -14'd1054,  -14'd829,  -14'd1185,  -14'd703,  
14'd519,  14'd119,  -14'd2233,  14'd456,  -14'd156,  -14'd664,  14'd2124,  -14'd1621,  14'd1008,  14'd438,  14'd633,  14'd1281,  14'd315,  -14'd478,  -14'd976,  14'd341,  
14'd194,  14'd816,  -14'd1101,  -14'd1667,  14'd1659,  -14'd914,  14'd757,  -14'd1129,  14'd795,  14'd769,  -14'd134,  14'd436,  -14'd322,  -14'd1296,  -14'd1838,  -14'd83,  
14'd1006,  14'd1681,  14'd263,  -14'd2442,  14'd2344,  -14'd411,  14'd767,  -14'd1233,  -14'd124,  14'd3074,  -14'd1643,  -14'd180,  -14'd1636,  14'd1423,  -14'd1198,  14'd628,  
-14'd1027,  14'd350,  14'd550,  14'd21,  14'd726,  -14'd617,  14'd1886,  -14'd1339,  14'd173,  -14'd1352,  -14'd1856,  -14'd322,  -14'd212,  14'd919,  14'd21,  -14'd995,  
14'd67,  -14'd160,  14'd1774,  -14'd762,  -14'd867,  14'd543,  14'd541,  -14'd1023,  14'd1355,  14'd710,  -14'd1308,  14'd366,  -14'd994,  14'd658,  14'd68,  -14'd208,  

-14'd2686,  -14'd885,  -14'd1358,  14'd594,  14'd308,  14'd97,  -14'd1600,  14'd674,  14'd634,  -14'd116,  -14'd1006,  -14'd448,  14'd405,  -14'd780,  -14'd315,  14'd970,  
14'd331,  -14'd1245,  14'd1321,  -14'd1004,  14'd405,  -14'd867,  14'd50,  14'd405,  -14'd31,  -14'd1220,  -14'd1352,  -14'd1287,  -14'd105,  14'd831,  -14'd868,  -14'd71,  
-14'd1416,  -14'd623,  14'd130,  14'd394,  -14'd650,  -14'd897,  -14'd42,  -14'd160,  -14'd1381,  14'd88,  -14'd640,  -14'd796,  -14'd382,  14'd3245,  14'd195,  -14'd2022,  
14'd804,  -14'd1047,  14'd1568,  -14'd248,  -14'd1208,  -14'd450,  -14'd97,  14'd359,  14'd69,  -14'd1011,  14'd291,  -14'd127,  -14'd1733,  -14'd72,  14'd435,  -14'd2106,  
14'd1487,  -14'd8,  -14'd440,  14'd1406,  -14'd808,  14'd1399,  -14'd817,  14'd545,  14'd642,  14'd778,  14'd326,  14'd27,  14'd1396,  -14'd1146,  14'd647,  14'd1240,  
-14'd523,  14'd763,  -14'd477,  14'd1060,  14'd853,  -14'd523,  -14'd1561,  -14'd1210,  -14'd1117,  14'd385,  -14'd239,  14'd271,  -14'd583,  14'd436,  14'd17,  -14'd372,  
14'd80,  -14'd1064,  -14'd20,  -14'd1013,  14'd947,  -14'd222,  14'd295,  14'd221,  -14'd277,  14'd464,  -14'd428,  14'd1220,  -14'd1965,  14'd549,  14'd330,  14'd44,  
14'd693,  14'd1314,  14'd1416,  14'd747,  14'd61,  14'd458,  -14'd1298,  14'd857,  14'd588,  14'd438,  14'd81,  -14'd484,  -14'd43,  14'd1880,  14'd515,  -14'd955,  
14'd14,  14'd217,  -14'd267,  14'd934,  -14'd1157,  14'd1259,  -14'd1207,  14'd1585,  -14'd1034,  -14'd338,  -14'd10,  -14'd1146,  14'd964,  -14'd89,  14'd93,  -14'd1071,  
14'd1520,  14'd527,  -14'd767,  14'd640,  14'd17,  14'd763,  -14'd1338,  -14'd484,  -14'd509,  14'd2347,  14'd723,  -14'd992,  14'd1432,  -14'd1158,  14'd779,  14'd1237,  
14'd183,  -14'd483,  14'd191,  14'd801,  -14'd1795,  14'd1076,  -14'd2083,  14'd877,  14'd809,  14'd27,  14'd1373,  14'd797,  14'd530,  -14'd366,  14'd213,  -14'd143,  
14'd490,  -14'd1773,  14'd282,  14'd570,  14'd1159,  14'd354,  14'd47,  14'd419,  14'd1430,  14'd69,  14'd954,  14'd1114,  14'd686,  -14'd520,  14'd893,  14'd127,  
-14'd695,  14'd591,  14'd1660,  14'd200,  -14'd673,  -14'd851,  14'd220,  -14'd449,  14'd1038,  14'd147,  14'd528,  14'd1766,  14'd72,  14'd1810,  14'd220,  -14'd476,  
-14'd1596,  -14'd61,  14'd1155,  14'd230,  -14'd401,  14'd0,  14'd1087,  -14'd122,  -14'd590,  14'd1266,  14'd1474,  14'd303,  -14'd248,  -14'd565,  14'd209,  -14'd1570,  
-14'd1678,  -14'd901,  14'd262,  14'd1729,  14'd178,  14'd81,  -14'd1382,  -14'd803,  14'd9,  14'd400,  14'd53,  -14'd170,  -14'd500,  -14'd878,  14'd409,  -14'd290,  
14'd886,  14'd533,  14'd409,  -14'd216,  -14'd192,  14'd263,  14'd1028,  14'd402,  14'd997,  14'd457,  14'd3057,  -14'd1146,  14'd1806,  -14'd209,  14'd240,  -14'd67,  
-14'd555,  14'd615,  14'd44,  14'd1027,  -14'd689,  14'd627,  14'd1256,  14'd989,  -14'd91,  14'd317,  14'd15,  14'd987,  -14'd132,  -14'd207,  14'd207,  -14'd986,  
14'd291,  -14'd352,  14'd125,  -14'd376,  -14'd480,  14'd440,  -14'd1143,  14'd12,  14'd1307,  -14'd478,  14'd796,  -14'd886,  14'd721,  14'd2852,  14'd349,  -14'd149,  
-14'd1188,  -14'd434,  14'd863,  -14'd93,  14'd358,  -14'd1256,  14'd162,  14'd479,  14'd283,  -14'd745,  14'd781,  -14'd663,  14'd374,  14'd350,  14'd967,  14'd1126,  
14'd837,  14'd1191,  14'd2516,  14'd495,  -14'd648,  14'd1040,  -14'd0,  -14'd7,  -14'd2,  14'd114,  14'd254,  14'd2071,  -14'd159,  -14'd71,  14'd251,  14'd431,  
14'd83,  14'd537,  -14'd1239,  -14'd637,  -14'd786,  -14'd1005,  14'd3108,  -14'd912,  14'd675,  -14'd1676,  14'd989,  -14'd604,  -14'd260,  -14'd233,  14'd206,  14'd859,  
14'd740,  14'd151,  14'd295,  -14'd544,  14'd373,  14'd764,  14'd1765,  14'd36,  14'd710,  14'd804,  -14'd238,  14'd770,  -14'd361,  14'd921,  -14'd537,  -14'd897,  
-14'd58,  -14'd411,  -14'd1085,  -14'd1184,  14'd688,  14'd51,  -14'd500,  14'd604,  -14'd187,  -14'd1097,  14'd436,  14'd115,  -14'd850,  14'd1818,  -14'd499,  14'd1304,  
-14'd2636,  -14'd215,  14'd750,  -14'd254,  -14'd643,  14'd41,  14'd538,  14'd856,  14'd690,  14'd168,  -14'd1487,  14'd1036,  -14'd234,  14'd96,  14'd1614,  14'd630,  
14'd2620,  14'd2045,  14'd1637,  -14'd1317,  14'd108,  14'd223,  -14'd1064,  -14'd345,  -14'd628,  -14'd113,  14'd1334,  14'd444,  14'd482,  -14'd395,  -14'd355,  14'd1240,  

14'd6,  14'd1133,  -14'd1469,  14'd889,  -14'd844,  14'd1196,  -14'd1663,  -14'd647,  -14'd18,  14'd761,  14'd1738,  14'd267,  14'd1843,  -14'd788,  -14'd91,  -14'd1006,  
14'd473,  -14'd566,  14'd19,  14'd492,  14'd411,  14'd1455,  -14'd598,  -14'd1471,  14'd622,  14'd226,  -14'd283,  14'd507,  14'd1160,  -14'd1940,  -14'd1016,  -14'd212,  
14'd1023,  -14'd582,  -14'd675,  -14'd340,  14'd1257,  14'd1329,  14'd647,  -14'd1196,  -14'd1215,  -14'd800,  14'd829,  14'd200,  14'd1293,  -14'd522,  -14'd1527,  -14'd1040,  
14'd1012,  14'd1808,  14'd447,  14'd868,  14'd1153,  14'd565,  -14'd500,  14'd322,  14'd978,  -14'd195,  14'd628,  -14'd347,  -14'd1318,  14'd1394,  14'd614,  14'd766,  
-14'd415,  14'd321,  14'd840,  14'd110,  -14'd1532,  -14'd120,  -14'd424,  -14'd365,  -14'd278,  -14'd9,  -14'd728,  -14'd794,  -14'd2726,  -14'd1863,  14'd1358,  -14'd714,  
14'd453,  14'd570,  -14'd2427,  14'd119,  -14'd761,  14'd102,  14'd680,  14'd498,  14'd950,  -14'd734,  14'd1581,  14'd518,  14'd752,  -14'd1225,  -14'd1424,  -14'd79,  
14'd206,  14'd589,  -14'd1086,  14'd573,  -14'd940,  -14'd504,  14'd469,  14'd614,  -14'd277,  14'd43,  14'd1041,  14'd1162,  14'd1672,  -14'd1473,  -14'd2267,  14'd671,  
14'd1182,  14'd1712,  -14'd405,  -14'd1006,  -14'd112,  -14'd295,  14'd1189,  -14'd1734,  14'd797,  -14'd1092,  14'd326,  14'd326,  14'd898,  14'd1638,  -14'd498,  14'd1837,  
-14'd115,  14'd1465,  14'd1277,  -14'd1687,  14'd1125,  14'd810,  14'd501,  14'd221,  -14'd227,  14'd248,  -14'd482,  -14'd830,  -14'd271,  14'd2164,  -14'd1066,  -14'd693,  
14'd328,  14'd941,  14'd954,  14'd493,  -14'd1189,  14'd303,  14'd1150,  14'd1175,  -14'd946,  -14'd15,  14'd420,  -14'd754,  -14'd2105,  -14'd238,  14'd127,  -14'd2242,  
-14'd618,  -14'd1412,  -14'd949,  -14'd1886,  -14'd346,  -14'd1897,  14'd929,  -14'd435,  -14'd541,  -14'd517,  14'd1329,  -14'd585,  -14'd1173,  -14'd722,  14'd806,  -14'd869,  
-14'd326,  -14'd1666,  -14'd916,  14'd320,  -14'd1582,  -14'd327,  -14'd1206,  -14'd1274,  14'd314,  14'd20,  14'd842,  14'd73,  -14'd750,  14'd356,  -14'd2464,  14'd898,  
-14'd10,  -14'd361,  -14'd1409,  -14'd1725,  14'd1413,  -14'd985,  14'd712,  -14'd981,  14'd739,  14'd1747,  14'd129,  -14'd646,  14'd509,  14'd891,  -14'd676,  -14'd689,  
14'd121,  14'd575,  14'd969,  -14'd1676,  14'd522,  -14'd836,  14'd583,  -14'd1295,  14'd814,  14'd124,  14'd224,  -14'd325,  14'd32,  14'd2092,  -14'd1032,  -14'd582,  
14'd2461,  14'd1204,  -14'd100,  14'd714,  -14'd723,  -14'd22,  14'd1144,  14'd650,  14'd940,  14'd493,  14'd1099,  -14'd687,  -14'd324,  -14'd1013,  -14'd131,  -14'd389,  
-14'd690,  -14'd445,  14'd337,  14'd713,  -14'd977,  -14'd447,  -14'd173,  -14'd1166,  -14'd153,  -14'd666,  -14'd236,  14'd433,  -14'd1155,  -14'd416,  -14'd41,  -14'd1291,  
14'd425,  -14'd1755,  -14'd1166,  -14'd1386,  14'd665,  -14'd1002,  -14'd1171,  -14'd1261,  14'd1002,  -14'd720,  14'd465,  14'd729,  14'd242,  -14'd390,  -14'd1023,  -14'd1199,  
-14'd72,  -14'd1080,  14'd121,  -14'd601,  14'd295,  -14'd1924,  14'd481,  -14'd1016,  14'd1223,  14'd276,  -14'd984,  14'd1521,  -14'd887,  -14'd683,  -14'd491,  -14'd692,  
14'd360,  -14'd1007,  14'd457,  -14'd39,  14'd449,  -14'd204,  -14'd834,  14'd235,  14'd1674,  14'd295,  -14'd1184,  -14'd977,  14'd307,  14'd1805,  14'd78,  -14'd1308,  
14'd135,  -14'd266,  -14'd2026,  -14'd946,  -14'd443,  14'd1272,  -14'd191,  14'd1063,  14'd2425,  14'd1090,  14'd338,  14'd776,  14'd738,  -14'd1938,  14'd1634,  -14'd909,  
14'd1014,  14'd0,  14'd795,  14'd846,  -14'd1983,  14'd415,  -14'd216,  -14'd313,  14'd48,  -14'd1991,  14'd634,  14'd210,  14'd522,  -14'd364,  -14'd108,  14'd95,  
14'd498,  -14'd1364,  -14'd1486,  14'd1485,  -14'd1495,  14'd913,  -14'd436,  14'd391,  14'd65,  -14'd107,  14'd1352,  14'd18,  14'd364,  -14'd98,  -14'd277,  14'd1332,  
14'd788,  14'd363,  14'd19,  14'd936,  -14'd1154,  14'd1585,  14'd165,  14'd371,  14'd310,  -14'd752,  14'd1639,  -14'd289,  14'd1734,  14'd260,  14'd802,  -14'd78,  
-14'd1434,  14'd484,  14'd897,  14'd682,  14'd1532,  14'd1073,  -14'd1041,  -14'd286,  -14'd187,  14'd2003,  14'd571,  -14'd403,  14'd604,  -14'd1923,  14'd590,  14'd1064,  
-14'd1334,  -14'd779,  14'd500,  14'd587,  -14'd120,  14'd1312,  14'd198,  14'd514,  14'd588,  14'd1632,  14'd1497,  14'd1280,  14'd785,  -14'd493,  14'd321,  14'd613,  

-14'd1082,  -14'd1111,  14'd281,  14'd873,  -14'd100,  14'd337,  -14'd220,  -14'd937,  14'd277,  14'd303,  14'd277,  -14'd123,  -14'd1191,  -14'd469,  14'd1118,  14'd194,  
14'd129,  14'd437,  14'd409,  -14'd553,  14'd288,  -14'd1200,  14'd392,  -14'd551,  -14'd462,  -14'd522,  -14'd8,  -14'd1321,  14'd390,  14'd667,  -14'd31,  -14'd752,  
14'd792,  -14'd432,  -14'd1137,  14'd314,  14'd675,  -14'd1732,  -14'd47,  14'd36,  -14'd141,  -14'd411,  -14'd418,  14'd275,  14'd637,  14'd1118,  14'd185,  -14'd561,  
14'd778,  -14'd331,  -14'd547,  14'd771,  -14'd974,  14'd1039,  -14'd861,  14'd90,  -14'd293,  14'd436,  -14'd696,  -14'd479,  -14'd1018,  14'd1057,  14'd582,  -14'd1079,  
14'd958,  14'd43,  14'd126,  -14'd807,  -14'd92,  -14'd223,  14'd30,  14'd1483,  14'd489,  -14'd1161,  -14'd737,  14'd378,  14'd7,  14'd602,  -14'd223,  -14'd1266,  
14'd34,  -14'd81,  14'd1278,  -14'd1014,  -14'd729,  14'd1470,  -14'd63,  -14'd456,  -14'd559,  14'd1028,  -14'd855,  14'd571,  14'd355,  -14'd1166,  -14'd438,  -14'd272,  
14'd739,  14'd819,  -14'd251,  -14'd428,  -14'd250,  -14'd977,  -14'd780,  -14'd573,  14'd1343,  -14'd1348,  -14'd478,  -14'd1027,  -14'd729,  -14'd1758,  14'd1231,  -14'd1670,  
14'd263,  14'd313,  -14'd210,  -14'd793,  -14'd772,  -14'd410,  -14'd261,  14'd19,  -14'd211,  -14'd955,  14'd911,  14'd772,  14'd792,  -14'd247,  14'd426,  14'd580,  
14'd648,  14'd967,  14'd375,  -14'd571,  -14'd150,  14'd108,  -14'd1513,  14'd810,  -14'd838,  -14'd846,  14'd412,  -14'd1707,  14'd417,  -14'd370,  -14'd732,  -14'd1676,  
-14'd257,  -14'd302,  14'd205,  14'd269,  -14'd754,  14'd285,  -14'd187,  -14'd118,  -14'd1120,  -14'd649,  -14'd901,  14'd989,  14'd307,  -14'd622,  14'd581,  -14'd1125,  
14'd772,  14'd272,  14'd419,  14'd463,  14'd297,  14'd299,  -14'd594,  14'd8,  -14'd212,  -14'd596,  -14'd241,  14'd86,  14'd223,  -14'd780,  -14'd385,  14'd63,  
14'd767,  -14'd574,  14'd770,  14'd1479,  -14'd581,  14'd112,  -14'd1298,  -14'd1256,  14'd278,  -14'd242,  -14'd351,  -14'd1219,  14'd1391,  -14'd55,  -14'd291,  -14'd452,  
14'd435,  14'd357,  -14'd687,  -14'd791,  14'd180,  -14'd1475,  14'd764,  -14'd1163,  14'd1089,  14'd1131,  14'd847,  -14'd775,  -14'd310,  -14'd557,  -14'd1518,  -14'd337,  
14'd205,  -14'd949,  14'd408,  14'd931,  -14'd615,  -14'd457,  -14'd160,  14'd529,  14'd1269,  -14'd763,  14'd276,  -14'd927,  14'd439,  14'd759,  14'd1372,  14'd546,  
14'd660,  -14'd1259,  14'd168,  14'd252,  -14'd459,  14'd52,  14'd794,  14'd534,  -14'd309,  -14'd636,  -14'd217,  -14'd354,  -14'd829,  14'd667,  14'd109,  -14'd571,  
-14'd298,  14'd100,  14'd1144,  -14'd486,  -14'd559,  -14'd962,  14'd216,  -14'd40,  14'd80,  14'd404,  -14'd421,  -14'd512,  -14'd531,  -14'd548,  -14'd96,  -14'd565,  
14'd496,  -14'd297,  -14'd658,  -14'd1072,  14'd358,  -14'd1003,  -14'd271,  14'd321,  -14'd769,  14'd555,  -14'd421,  14'd405,  -14'd1206,  14'd877,  -14'd286,  -14'd235,  
-14'd188,  -14'd682,  -14'd117,  -14'd112,  -14'd41,  14'd213,  -14'd833,  -14'd934,  14'd181,  -14'd764,  -14'd32,  -14'd931,  14'd3,  -14'd222,  -14'd979,  14'd310,  
14'd501,  -14'd279,  -14'd580,  -14'd727,  -14'd1258,  14'd794,  -14'd9,  -14'd453,  -14'd156,  14'd71,  14'd305,  -14'd1177,  -14'd320,  -14'd1776,  -14'd164,  -14'd224,  
14'd1549,  -14'd937,  -14'd543,  -14'd516,  -14'd523,  -14'd112,  -14'd114,  -14'd280,  14'd497,  -14'd73,  14'd59,  14'd173,  14'd1044,  14'd749,  -14'd63,  -14'd1644,  
14'd354,  -14'd90,  -14'd153,  -14'd1416,  -14'd389,  14'd1260,  -14'd90,  -14'd229,  -14'd20,  14'd1123,  -14'd1220,  -14'd261,  -14'd865,  14'd523,  14'd668,  -14'd371,  
-14'd277,  -14'd1743,  -14'd1034,  -14'd89,  -14'd659,  -14'd431,  -14'd443,  14'd884,  14'd656,  -14'd36,  -14'd1018,  -14'd712,  -14'd1321,  -14'd1484,  -14'd7,  14'd913,  
-14'd480,  -14'd291,  14'd589,  14'd119,  14'd305,  14'd600,  -14'd353,  -14'd1167,  14'd176,  -14'd482,  -14'd1073,  -14'd1663,  -14'd827,  14'd1034,  -14'd907,  14'd21,  
14'd501,  14'd485,  -14'd620,  -14'd1193,  14'd1284,  -14'd1199,  -14'd633,  -14'd828,  14'd842,  14'd1081,  -14'd722,  14'd150,  -14'd425,  -14'd279,  -14'd792,  -14'd89,  
14'd604,  14'd111,  -14'd189,  -14'd87,  -14'd347,  -14'd218,  -14'd796,  -14'd967,  -14'd207,  14'd309,  -14'd120,  -14'd403,  -14'd779,  14'd1003,  -14'd978,  -14'd191,  

14'd522,  -14'd151,  -14'd1534,  -14'd1211,  -14'd922,  -14'd2574,  14'd2543,  -14'd1980,  14'd215,  -14'd2308,  -14'd2014,  -14'd155,  -14'd1199,  14'd906,  -14'd1864,  -14'd1653,  
-14'd141,  14'd846,  -14'd1727,  -14'd312,  -14'd352,  -14'd1449,  -14'd28,  14'd55,  14'd55,  14'd1068,  -14'd2081,  -14'd167,  -14'd1518,  -14'd1040,  -14'd283,  -14'd1694,  
14'd1621,  14'd1017,  -14'd1557,  -14'd115,  -14'd323,  14'd1597,  -14'd2000,  14'd1172,  -14'd247,  14'd308,  14'd330,  14'd536,  14'd154,  -14'd3036,  14'd1109,  14'd955,  
14'd196,  -14'd725,  -14'd368,  14'd424,  14'd575,  14'd457,  -14'd11,  -14'd304,  14'd936,  14'd683,  14'd803,  14'd1132,  14'd226,  -14'd1563,  14'd702,  14'd316,  
-14'd2334,  14'd949,  14'd109,  -14'd749,  -14'd162,  14'd425,  14'd4,  -14'd858,  -14'd282,  -14'd557,  14'd731,  14'd401,  -14'd853,  14'd240,  14'd365,  14'd1034,  
-14'd350,  -14'd41,  -14'd1269,  14'd80,  -14'd1516,  -14'd382,  14'd28,  14'd181,  -14'd840,  14'd594,  -14'd869,  -14'd62,  14'd254,  -14'd188,  -14'd885,  -14'd1610,  
14'd1320,  14'd600,  14'd643,  -14'd621,  14'd461,  -14'd185,  -14'd216,  14'd918,  14'd252,  -14'd380,  -14'd1319,  -14'd594,  -14'd938,  -14'd121,  14'd496,  -14'd75,  
14'd471,  -14'd329,  -14'd163,  -14'd838,  -14'd1332,  -14'd430,  14'd84,  14'd1768,  14'd451,  14'd139,  -14'd295,  14'd230,  -14'd939,  -14'd2680,  14'd1799,  -14'd510,  
14'd1031,  -14'd1002,  14'd80,  14'd174,  -14'd249,  14'd647,  14'd277,  14'd135,  -14'd247,  -14'd704,  -14'd893,  -14'd1038,  14'd346,  14'd663,  -14'd150,  14'd191,  
-14'd1744,  -14'd531,  -14'd709,  14'd552,  -14'd509,  14'd302,  14'd1434,  14'd818,  14'd1234,  -14'd1263,  14'd1638,  14'd703,  -14'd86,  14'd1347,  -14'd423,  -14'd625,  
14'd1233,  14'd631,  14'd1481,  -14'd97,  14'd1181,  -14'd149,  14'd190,  -14'd501,  -14'd457,  -14'd21,  -14'd2954,  14'd383,  -14'd336,  14'd1393,  14'd305,  14'd246,  
-14'd85,  -14'd657,  14'd1592,  -14'd455,  14'd910,  14'd405,  -14'd1400,  14'd647,  14'd12,  14'd179,  -14'd1689,  14'd532,  14'd364,  14'd716,  14'd65,  -14'd1680,  
14'd225,  -14'd168,  14'd1412,  14'd851,  -14'd531,  -14'd5,  14'd563,  -14'd848,  14'd66,  -14'd656,  14'd726,  -14'd304,  -14'd998,  -14'd710,  14'd367,  14'd238,  
14'd677,  14'd1140,  14'd396,  -14'd1539,  14'd372,  -14'd870,  -14'd244,  -14'd317,  14'd692,  14'd284,  14'd949,  -14'd1218,  -14'd212,  14'd1338,  -14'd945,  14'd507,  
-14'd453,  14'd4,  14'd765,  -14'd732,  14'd37,  14'd315,  14'd45,  14'd860,  14'd455,  -14'd1739,  14'd782,  -14'd539,  14'd316,  14'd2165,  14'd1426,  -14'd143,  
14'd121,  14'd50,  14'd899,  14'd520,  -14'd471,  -14'd164,  -14'd2347,  14'd234,  -14'd1462,  14'd391,  -14'd1748,  14'd74,  14'd69,  14'd716,  -14'd216,  -14'd13,  
-14'd295,  -14'd91,  14'd1044,  14'd679,  -14'd95,  -14'd187,  14'd67,  -14'd183,  -14'd326,  -14'd560,  -14'd981,  14'd200,  -14'd128,  14'd513,  -14'd13,  -14'd778,  
-14'd588,  14'd2301,  14'd1134,  -14'd1658,  14'd1215,  -14'd854,  14'd526,  -14'd495,  -14'd611,  14'd508,  -14'd34,  14'd546,  -14'd336,  -14'd153,  14'd1427,  -14'd365,  
-14'd162,  14'd181,  14'd1296,  -14'd16,  -14'd201,  -14'd475,  14'd1032,  -14'd1450,  14'd277,  -14'd1340,  -14'd1288,  14'd1302,  14'd254,  14'd1218,  -14'd1669,  -14'd177,  
14'd705,  14'd1362,  -14'd744,  -14'd1179,  -14'd1269,  -14'd33,  -14'd587,  14'd619,  -14'd744,  -14'd1938,  -14'd914,  -14'd1044,  14'd293,  14'd867,  -14'd1937,  -14'd2332,  
-14'd1339,  14'd148,  14'd833,  14'd869,  14'd2021,  14'd715,  -14'd1130,  14'd72,  -14'd609,  14'd408,  14'd798,  -14'd5,  -14'd284,  -14'd74,  -14'd263,  -14'd651,  
14'd285,  14'd115,  -14'd194,  -14'd1045,  14'd209,  -14'd443,  -14'd1551,  -14'd416,  -14'd719,  -14'd1509,  14'd594,  14'd509,  14'd514,  -14'd403,  14'd61,  14'd916,  
14'd1603,  -14'd1447,  -14'd361,  14'd1153,  -14'd297,  -14'd202,  -14'd685,  -14'd668,  14'd1471,  14'd541,  -14'd363,  14'd659,  -14'd66,  -14'd1133,  -14'd322,  14'd37,  
14'd1831,  -14'd414,  14'd1010,  14'd486,  -14'd418,  -14'd590,  14'd385,  14'd686,  14'd600,  14'd765,  14'd98,  14'd1591,  14'd361,  14'd617,  -14'd1381,  14'd166,  
14'd373,  -14'd954,  -14'd1436,  -14'd1046,  -14'd1055,  -14'd1311,  -14'd294,  14'd923,  14'd1869,  -14'd2107,  -14'd1065,  -14'd2043,  14'd101,  14'd830,  -14'd402,  -14'd284,  

14'd244,  -14'd549,  -14'd213,  14'd24,  14'd68,  14'd1046,  -14'd2316,  14'd34,  14'd450,  -14'd182,  14'd788,  -14'd1033,  -14'd191,  -14'd2096,  14'd119,  -14'd488,  
-14'd112,  14'd531,  -14'd314,  14'd886,  14'd24,  -14'd557,  -14'd607,  -14'd110,  14'd1859,  14'd552,  -14'd1119,  -14'd1662,  14'd774,  -14'd343,  -14'd385,  14'd2548,  
-14'd274,  -14'd1133,  -14'd273,  -14'd1415,  14'd1535,  14'd137,  -14'd205,  14'd1409,  14'd208,  14'd109,  -14'd1852,  14'd600,  14'd610,  -14'd6,  -14'd330,  14'd575,  
-14'd1445,  -14'd1834,  -14'd864,  -14'd664,  14'd894,  -14'd885,  14'd277,  -14'd333,  -14'd227,  -14'd1902,  -14'd782,  -14'd933,  -14'd654,  14'd2308,  -14'd1096,  14'd634,  
-14'd699,  -14'd294,  14'd761,  -14'd851,  14'd873,  -14'd27,  -14'd797,  14'd108,  -14'd301,  -14'd283,  -14'd902,  14'd1330,  -14'd1334,  14'd673,  14'd425,  -14'd1895,  
14'd319,  14'd537,  -14'd1210,  -14'd644,  14'd1735,  -14'd1112,  -14'd762,  14'd989,  -14'd113,  -14'd1060,  -14'd190,  -14'd149,  14'd96,  -14'd2294,  14'd673,  -14'd402,  
-14'd182,  14'd51,  -14'd168,  -14'd1529,  14'd125,  -14'd518,  14'd680,  -14'd63,  -14'd6,  14'd925,  -14'd830,  14'd994,  -14'd760,  14'd204,  14'd748,  14'd443,  
14'd1646,  -14'd813,  14'd719,  -14'd463,  14'd653,  14'd410,  14'd515,  14'd1363,  -14'd143,  14'd1397,  -14'd248,  14'd1866,  -14'd753,  14'd1419,  14'd1112,  14'd895,  
14'd2415,  -14'd1365,  14'd1450,  14'd507,  14'd21,  14'd1147,  14'd421,  14'd1261,  -14'd122,  -14'd574,  14'd356,  14'd1133,  -14'd210,  14'd1959,  14'd591,  14'd1101,  
14'd1766,  14'd1136,  -14'd372,  14'd32,  14'd1157,  14'd905,  -14'd210,  -14'd432,  14'd104,  -14'd1830,  -14'd1535,  -14'd1157,  14'd1163,  14'd1394,  -14'd482,  -14'd300,  
-14'd159,  -14'd273,  -14'd57,  14'd470,  14'd531,  14'd734,  -14'd488,  14'd635,  14'd1180,  -14'd68,  14'd175,  -14'd1254,  14'd393,  -14'd1033,  14'd683,  14'd400,  
14'd460,  -14'd855,  -14'd897,  -14'd629,  -14'd1097,  14'd707,  -14'd366,  14'd974,  14'd1075,  14'd638,  14'd22,  14'd217,  14'd1807,  14'd901,  -14'd43,  -14'd20,  
-14'd66,  -14'd626,  -14'd1763,  14'd1774,  -14'd1091,  -14'd540,  -14'd104,  14'd417,  -14'd190,  14'd982,  14'd1515,  14'd1145,  14'd783,  -14'd1426,  14'd495,  14'd1359,  
-14'd136,  -14'd2251,  14'd1797,  14'd736,  14'd477,  14'd336,  14'd457,  14'd1625,  -14'd782,  14'd3,  14'd579,  14'd1018,  14'd1622,  -14'd1577,  14'd345,  -14'd95,  
-14'd249,  -14'd772,  -14'd1145,  -14'd331,  -14'd1048,  -14'd371,  14'd1265,  14'd1386,  -14'd333,  14'd436,  -14'd81,  -14'd1243,  14'd1655,  -14'd181,  -14'd108,  14'd1445,  
-14'd207,  -14'd1030,  14'd1352,  -14'd142,  14'd1168,  -14'd71,  -14'd1394,  14'd587,  14'd210,  -14'd50,  -14'd30,  -14'd20,  14'd599,  -14'd922,  -14'd90,  -14'd673,  
-14'd1006,  14'd295,  14'd101,  14'd301,  14'd477,  -14'd718,  -14'd1050,  14'd622,  14'd663,  -14'd511,  -14'd747,  14'd595,  14'd474,  14'd169,  -14'd18,  14'd1080,  
-14'd615,  -14'd711,  -14'd1032,  14'd165,  -14'd45,  -14'd807,  14'd26,  -14'd916,  -14'd978,  -14'd260,  -14'd310,  14'd226,  -14'd1087,  -14'd899,  -14'd739,  14'd146,  
14'd1000,  14'd1357,  14'd409,  -14'd718,  -14'd2112,  14'd1324,  -14'd843,  14'd53,  14'd492,  14'd502,  14'd946,  14'd398,  -14'd402,  -14'd234,  14'd423,  14'd342,  
-14'd676,  14'd269,  -14'd524,  -14'd38,  14'd1515,  -14'd618,  14'd367,  14'd1460,  14'd494,  -14'd1050,  14'd210,  14'd990,  -14'd423,  14'd542,  14'd875,  -14'd298,  
-14'd256,  14'd326,  -14'd620,  14'd1288,  14'd733,  14'd692,  -14'd588,  -14'd563,  -14'd107,  -14'd628,  -14'd252,  14'd1515,  14'd349,  14'd321,  -14'd550,  -14'd616,  
14'd364,  14'd462,  -14'd1450,  14'd261,  -14'd1117,  -14'd891,  -14'd1768,  -14'd1221,  14'd328,  14'd776,  14'd479,  -14'd24,  -14'd825,  14'd472,  14'd582,  14'd507,  
-14'd71,  -14'd582,  -14'd344,  -14'd1621,  14'd598,  -14'd1019,  14'd896,  14'd890,  14'd645,  14'd1073,  -14'd750,  14'd528,  -14'd802,  14'd1213,  14'd643,  -14'd384,  
14'd340,  -14'd933,  14'd1917,  -14'd586,  14'd341,  14'd336,  14'd1057,  -14'd549,  14'd1713,  -14'd727,  -14'd437,  14'd861,  -14'd811,  14'd315,  14'd603,  14'd167,  
14'd101,  -14'd380,  14'd804,  -14'd456,  14'd387,  -14'd618,  14'd1575,  14'd1250,  -14'd832,  -14'd2475,  -14'd227,  14'd989,  14'd185,  -14'd21,  -14'd484,  14'd518,  

14'd1551,  14'd701,  -14'd1198,  -14'd574,  -14'd708,  14'd1745,  -14'd808,  14'd479,  -14'd304,  14'd91,  14'd572,  14'd506,  14'd299,  -14'd1519,  14'd1274,  14'd491,  
-14'd570,  14'd558,  -14'd929,  -14'd821,  -14'd691,  14'd662,  14'd646,  14'd1779,  -14'd167,  14'd736,  14'd622,  14'd90,  -14'd278,  -14'd1250,  14'd1354,  14'd586,  
14'd196,  14'd1271,  -14'd1473,  14'd456,  14'd641,  14'd488,  -14'd106,  -14'd1150,  -14'd676,  14'd170,  14'd107,  14'd333,  -14'd1240,  14'd1864,  14'd334,  14'd717,  
14'd38,  14'd262,  14'd621,  -14'd1385,  -14'd319,  14'd446,  14'd432,  -14'd1273,  14'd486,  14'd898,  -14'd818,  -14'd245,  -14'd67,  14'd959,  -14'd606,  -14'd812,  
-14'd500,  -14'd156,  -14'd1451,  -14'd262,  14'd1562,  14'd323,  -14'd701,  -14'd1315,  -14'd1531,  -14'd1121,  -14'd221,  -14'd456,  -14'd1733,  14'd1062,  14'd832,  14'd1109,  
14'd957,  -14'd675,  -14'd112,  14'd608,  14'd106,  -14'd881,  14'd713,  14'd646,  -14'd527,  14'd1448,  14'd102,  -14'd62,  14'd673,  -14'd382,  -14'd360,  14'd1139,  
14'd553,  14'd1059,  -14'd298,  14'd713,  14'd830,  -14'd36,  14'd661,  -14'd1332,  -14'd26,  14'd1486,  -14'd1303,  -14'd964,  14'd122,  14'd227,  -14'd221,  14'd1537,  
-14'd295,  14'd84,  -14'd739,  -14'd595,  14'd57,  -14'd1229,  -14'd1212,  14'd671,  -14'd1218,  14'd690,  14'd1296,  14'd719,  14'd844,  -14'd787,  14'd129,  14'd1082,  
14'd907,  -14'd1330,  14'd249,  14'd353,  -14'd371,  -14'd420,  -14'd682,  -14'd1119,  14'd197,  -14'd464,  -14'd280,  14'd171,  -14'd642,  14'd434,  -14'd1167,  14'd1119,  
14'd1951,  14'd2122,  14'd420,  -14'd1015,  -14'd165,  14'd386,  14'd584,  -14'd347,  14'd423,  -14'd594,  -14'd384,  14'd1579,  14'd899,  -14'd782,  -14'd1434,  -14'd1299,  
-14'd958,  14'd1251,  -14'd538,  -14'd418,  14'd437,  -14'd262,  -14'd401,  14'd447,  14'd171,  14'd1297,  14'd899,  14'd83,  14'd161,  -14'd115,  -14'd1091,  -14'd211,  
14'd1132,  14'd934,  14'd843,  -14'd72,  -14'd233,  14'd800,  -14'd943,  14'd725,  14'd474,  14'd368,  -14'd114,  14'd73,  -14'd242,  -14'd597,  -14'd300,  14'd857,  
14'd1411,  14'd760,  14'd625,  14'd232,  -14'd684,  14'd1753,  14'd668,  14'd288,  14'd1293,  -14'd210,  14'd1147,  14'd682,  -14'd711,  -14'd1436,  -14'd378,  14'd155,  
14'd1230,  -14'd2057,  14'd307,  -14'd206,  14'd704,  14'd421,  14'd341,  -14'd554,  14'd1255,  14'd912,  14'd144,  -14'd465,  -14'd403,  14'd307,  14'd1426,  14'd635,  
14'd609,  14'd247,  -14'd1807,  14'd1081,  -14'd114,  14'd895,  -14'd40,  -14'd567,  14'd357,  14'd1125,  14'd71,  -14'd155,  14'd774,  -14'd244,  -14'd130,  14'd950,  
14'd492,  -14'd204,  -14'd429,  -14'd423,  -14'd1057,  14'd196,  -14'd348,  -14'd1013,  14'd1086,  -14'd708,  -14'd1741,  14'd392,  14'd294,  14'd1050,  14'd240,  -14'd924,  
14'd1251,  14'd699,  14'd804,  14'd1324,  14'd253,  14'd468,  14'd108,  -14'd473,  14'd815,  14'd30,  -14'd225,  -14'd158,  14'd402,  14'd1718,  14'd209,  -14'd94,  
-14'd1153,  14'd475,  -14'd404,  14'd787,  -14'd806,  14'd361,  14'd180,  -14'd1077,  14'd1721,  14'd784,  -14'd311,  -14'd351,  14'd308,  -14'd2206,  -14'd384,  14'd173,  
-14'd749,  -14'd469,  14'd171,  14'd188,  14'd133,  14'd710,  14'd433,  14'd412,  -14'd755,  14'd403,  14'd1339,  -14'd686,  14'd377,  -14'd1454,  14'd417,  -14'd1349,  
-14'd1735,  -14'd3,  -14'd640,  14'd485,  14'd356,  14'd197,  -14'd491,  -14'd561,  -14'd366,  14'd507,  14'd359,  14'd539,  14'd535,  14'd27,  -14'd118,  14'd417,  
14'd1114,  -14'd284,  14'd1622,  14'd929,  -14'd849,  14'd826,  -14'd33,  14'd1418,  -14'd36,  14'd73,  -14'd1395,  14'd809,  14'd403,  14'd1502,  14'd620,  14'd42,  
14'd866,  14'd851,  14'd227,  14'd577,  14'd856,  -14'd720,  -14'd1630,  14'd2143,  -14'd201,  -14'd743,  -14'd1002,  -14'd59,  14'd1341,  14'd1127,  14'd140,  14'd15,  
-14'd1764,  -14'd584,  14'd89,  14'd564,  14'd1059,  14'd446,  14'd350,  14'd44,  -14'd2228,  -14'd3488,  14'd355,  14'd295,  14'd833,  -14'd1389,  14'd382,  -14'd754,  
-14'd1398,  14'd490,  -14'd1462,  -14'd354,  -14'd877,  -14'd11,  -14'd365,  14'd350,  14'd770,  -14'd1604,  14'd112,  14'd817,  -14'd379,  -14'd43,  14'd1027,  -14'd1042,  
-14'd681,  14'd719,  14'd476,  14'd790,  -14'd369,  -14'd212,  14'd650,  -14'd196,  14'd46,  -14'd1043,  14'd711,  14'd1082,  14'd466,  -14'd379,  -14'd251,  14'd76,  

14'd904,  14'd796,  14'd339,  14'd597,  -14'd2136,  14'd674,  14'd2455,  -14'd57,  14'd371,  -14'd1041,  -14'd1559,  14'd1155,  -14'd1941,  14'd184,  -14'd900,  14'd178,  
14'd238,  14'd161,  -14'd871,  -14'd1408,  -14'd868,  14'd653,  -14'd934,  -14'd1062,  14'd756,  14'd263,  14'd2010,  -14'd321,  -14'd1260,  14'd1203,  -14'd1042,  -14'd626,  
14'd420,  14'd266,  -14'd2174,  -14'd560,  14'd870,  14'd311,  -14'd946,  -14'd963,  -14'd698,  14'd763,  14'd379,  -14'd803,  -14'd847,  14'd1114,  -14'd862,  14'd1078,  
-14'd749,  14'd716,  14'd12,  14'd768,  14'd985,  -14'd366,  -14'd610,  -14'd434,  14'd481,  14'd497,  -14'd124,  -14'd228,  14'd187,  14'd102,  -14'd316,  -14'd435,  
14'd690,  14'd2461,  14'd681,  -14'd695,  14'd398,  14'd869,  -14'd364,  14'd1067,  -14'd675,  14'd258,  14'd387,  14'd643,  14'd1194,  14'd378,  14'd807,  14'd1073,  
14'd472,  -14'd321,  14'd455,  -14'd181,  14'd128,  14'd851,  -14'd505,  -14'd47,  -14'd407,  14'd635,  -14'd984,  14'd742,  -14'd121,  14'd2757,  -14'd545,  14'd534,  
14'd770,  -14'd311,  14'd562,  14'd618,  -14'd1127,  14'd164,  -14'd309,  14'd985,  14'd261,  14'd368,  -14'd839,  -14'd1341,  14'd1586,  14'd1376,  14'd1663,  -14'd76,  
-14'd1891,  -14'd1072,  14'd216,  -14'd1427,  -14'd596,  -14'd912,  -14'd520,  -14'd171,  14'd857,  14'd74,  14'd1041,  -14'd5,  -14'd903,  -14'd467,  14'd237,  -14'd596,  
-14'd2014,  -14'd758,  -14'd223,  -14'd858,  -14'd422,  14'd1564,  -14'd1214,  14'd743,  -14'd17,  -14'd127,  -14'd558,  14'd1006,  -14'd189,  -14'd280,  14'd580,  -14'd699,  
-14'd554,  14'd1145,  -14'd964,  -14'd219,  14'd714,  14'd481,  14'd560,  14'd391,  14'd870,  14'd928,  -14'd833,  -14'd878,  -14'd626,  14'd292,  -14'd250,  14'd188,  
14'd893,  14'd421,  -14'd269,  14'd1786,  14'd408,  14'd2732,  -14'd2283,  14'd1368,  -14'd1494,  14'd982,  -14'd871,  14'd1020,  14'd908,  14'd596,  14'd896,  14'd978,  
-14'd794,  14'd2039,  14'd580,  14'd912,  14'd1082,  -14'd636,  -14'd1874,  14'd1284,  14'd89,  -14'd1014,  14'd2092,  14'd1388,  -14'd804,  14'd373,  14'd57,  14'd1640,  
-14'd939,  -14'd631,  14'd488,  14'd885,  14'd141,  14'd702,  -14'd712,  14'd1558,  14'd1456,  -14'd2459,  14'd526,  -14'd324,  14'd382,  -14'd17,  14'd266,  -14'd67,  
-14'd333,  14'd37,  -14'd1304,  14'd161,  -14'd1505,  14'd18,  -14'd192,  -14'd60,  14'd645,  14'd81,  14'd33,  14'd354,  14'd240,  -14'd178,  -14'd1162,  14'd854,  
14'd342,  14'd81,  -14'd1248,  -14'd79,  14'd171,  14'd106,  -14'd1558,  14'd333,  -14'd806,  14'd188,  -14'd107,  -14'd230,  14'd457,  14'd111,  14'd88,  14'd783,  
14'd1455,  14'd1170,  -14'd291,  -14'd228,  14'd1526,  -14'd217,  -14'd1451,  14'd1053,  -14'd552,  -14'd226,  -14'd1195,  14'd1037,  14'd800,  14'd1128,  -14'd74,  14'd952,  
14'd299,  14'd1681,  14'd1538,  -14'd544,  14'd1166,  14'd1324,  14'd673,  -14'd640,  -14'd718,  14'd627,  -14'd90,  -14'd321,  -14'd1497,  14'd457,  14'd187,  14'd734,  
14'd142,  14'd376,  14'd187,  -14'd90,  14'd341,  14'd216,  14'd847,  -14'd608,  14'd2158,  -14'd65,  -14'd649,  -14'd342,  -14'd1030,  -14'd923,  -14'd600,  14'd750,  
-14'd1406,  14'd1185,  -14'd747,  -14'd623,  14'd887,  -14'd516,  14'd310,  14'd410,  -14'd692,  14'd353,  14'd96,  -14'd161,  -14'd1207,  14'd726,  -14'd418,  -14'd536,  
-14'd654,  -14'd1194,  14'd887,  -14'd297,  14'd402,  -14'd354,  14'd0,  -14'd930,  -14'd1664,  -14'd26,  14'd780,  14'd182,  -14'd856,  14'd49,  -14'd497,  -14'd5,  
14'd1619,  -14'd304,  14'd168,  14'd235,  -14'd61,  -14'd734,  14'd612,  14'd611,  14'd1203,  -14'd842,  -14'd1034,  14'd85,  14'd406,  14'd117,  14'd113,  -14'd145,  
-14'd1093,  -14'd617,  14'd0,  14'd94,  14'd65,  -14'd477,  -14'd1253,  14'd358,  -14'd273,  14'd828,  -14'd10,  -14'd826,  -14'd353,  -14'd42,  -14'd217,  -14'd20,  
-14'd597,  -14'd544,  14'd624,  14'd233,  -14'd729,  -14'd617,  -14'd1329,  14'd406,  -14'd212,  14'd411,  -14'd864,  -14'd183,  -14'd356,  -14'd560,  14'd692,  14'd420,  
-14'd1240,  14'd512,  -14'd269,  14'd1446,  -14'd237,  14'd792,  -14'd287,  -14'd303,  -14'd365,  -14'd864,  14'd28,  14'd986,  -14'd69,  14'd1585,  14'd205,  -14'd479,  
-14'd814,  -14'd967,  -14'd263,  14'd933,  -14'd779,  -14'd735,  -14'd6,  -14'd308,  14'd163,  -14'd1668,  -14'd832,  14'd591,  14'd350,  -14'd427,  14'd230,  14'd1473,  

-14'd343,  14'd73,  14'd34,  -14'd110,  14'd594,  -14'd349,  -14'd1549,  14'd1162,  -14'd94,  14'd377,  -14'd1938,  -14'd880,  14'd992,  -14'd25,  -14'd1598,  -14'd119,  
-14'd1332,  14'd533,  14'd1460,  14'd674,  14'd1421,  -14'd65,  -14'd1742,  -14'd900,  -14'd387,  14'd1032,  -14'd1124,  14'd537,  14'd596,  14'd1354,  14'd1219,  14'd1497,  
14'd143,  -14'd1061,  14'd513,  -14'd871,  14'd134,  -14'd875,  -14'd153,  14'd230,  14'd76,  -14'd607,  14'd141,  14'd1292,  -14'd493,  14'd1564,  14'd1097,  14'd1268,  
14'd116,  -14'd454,  14'd1093,  14'd573,  -14'd39,  14'd414,  14'd816,  14'd781,  -14'd233,  -14'd278,  14'd154,  14'd1004,  -14'd892,  14'd2088,  14'd1305,  -14'd244,  
14'd1230,  -14'd928,  14'd63,  -14'd447,  -14'd845,  -14'd672,  14'd1233,  -14'd691,  14'd1006,  -14'd38,  -14'd241,  14'd536,  -14'd844,  14'd457,  14'd601,  -14'd674,  
-14'd504,  -14'd902,  14'd449,  -14'd112,  14'd532,  14'd491,  -14'd1537,  14'd1034,  -14'd1539,  14'd307,  -14'd1057,  -14'd279,  -14'd445,  14'd850,  14'd236,  -14'd1189,  
14'd858,  14'd865,  14'd760,  14'd1499,  -14'd172,  14'd876,  14'd379,  -14'd292,  14'd473,  14'd16,  14'd885,  14'd1714,  -14'd709,  14'd5,  14'd722,  -14'd1309,  
-14'd394,  14'd992,  14'd1333,  14'd706,  14'd340,  14'd461,  14'd639,  14'd1427,  14'd1072,  14'd94,  14'd197,  -14'd435,  14'd57,  14'd2114,  14'd845,  -14'd1430,  
-14'd860,  14'd605,  14'd472,  14'd346,  -14'd543,  14'd316,  14'd472,  14'd623,  -14'd354,  -14'd1946,  14'd1035,  14'd794,  -14'd1473,  14'd160,  14'd513,  -14'd109,  
14'd730,  14'd922,  14'd44,  -14'd968,  14'd736,  14'd284,  14'd561,  -14'd678,  14'd833,  -14'd1325,  -14'd108,  -14'd667,  14'd124,  -14'd1655,  14'd587,  14'd887,  
14'd1285,  14'd11,  -14'd377,  -14'd379,  14'd286,  -14'd971,  -14'd263,  -14'd352,  14'd1441,  14'd258,  14'd2546,  -14'd680,  -14'd741,  14'd993,  14'd231,  -14'd99,  
14'd129,  14'd1081,  14'd356,  -14'd606,  -14'd1052,  14'd769,  14'd193,  14'd1466,  -14'd664,  14'd296,  14'd599,  -14'd109,  14'd254,  14'd117,  14'd221,  14'd1273,  
14'd400,  14'd859,  14'd649,  14'd599,  14'd358,  -14'd356,  14'd267,  14'd895,  -14'd607,  14'd192,  14'd20,  14'd785,  14'd367,  14'd1415,  -14'd200,  -14'd502,  
-14'd1087,  14'd285,  14'd967,  -14'd51,  -14'd21,  14'd81,  14'd1269,  14'd77,  -14'd426,  -14'd453,  14'd1370,  14'd371,  -14'd684,  -14'd694,  -14'd478,  -14'd1857,  
14'd670,  14'd17,  -14'd500,  14'd597,  14'd617,  14'd381,  14'd468,  14'd204,  -14'd72,  -14'd2835,  -14'd862,  -14'd1306,  -14'd550,  14'd100,  14'd476,  -14'd1365,  
-14'd151,  14'd855,  -14'd343,  -14'd398,  14'd2306,  -14'd1010,  -14'd1438,  14'd108,  14'd1239,  -14'd778,  14'd402,  -14'd292,  14'd334,  14'd98,  -14'd1709,  14'd154,  
-14'd449,  -14'd1263,  -14'd287,  14'd575,  -14'd54,  -14'd72,  14'd1074,  -14'd314,  -14'd425,  -14'd391,  14'd569,  14'd430,  -14'd47,  14'd503,  -14'd874,  14'd702,  
14'd1159,  -14'd343,  -14'd104,  14'd273,  -14'd465,  14'd1799,  -14'd231,  -14'd1186,  14'd443,  14'd63,  14'd382,  -14'd1218,  14'd692,  14'd811,  14'd402,  -14'd245,  
-14'd55,  -14'd973,  -14'd48,  14'd348,  14'd924,  -14'd1637,  -14'd1029,  -14'd4,  14'd2118,  14'd264,  14'd542,  -14'd521,  -14'd954,  14'd123,  14'd13,  14'd1034,  
14'd1152,  -14'd217,  14'd325,  -14'd799,  -14'd626,  -14'd672,  -14'd756,  -14'd84,  -14'd39,  14'd510,  -14'd943,  14'd334,  14'd470,  -14'd577,  -14'd530,  -14'd108,  
-14'd1163,  -14'd700,  -14'd1732,  -14'd293,  -14'd817,  14'd77,  -14'd101,  14'd316,  14'd816,  -14'd765,  14'd2035,  -14'd32,  -14'd423,  14'd312,  14'd140,  14'd367,  
-14'd177,  14'd661,  -14'd1353,  14'd18,  -14'd501,  14'd760,  14'd865,  -14'd2043,  14'd1556,  -14'd1194,  14'd562,  14'd1670,  -14'd1243,  14'd422,  14'd34,  14'd467,  
-14'd258,  14'd1003,  14'd393,  -14'd1506,  -14'd66,  -14'd75,  14'd1064,  -14'd708,  14'd852,  14'd1229,  14'd454,  -14'd61,  14'd230,  14'd1706,  14'd215,  14'd1473,  
14'd564,  -14'd51,  14'd1341,  14'd1105,  -14'd286,  -14'd941,  -14'd443,  -14'd419,  -14'd960,  14'd548,  -14'd1032,  -14'd706,  -14'd1560,  14'd492,  14'd754,  -14'd509,  
14'd1663,  14'd1481,  14'd1608,  -14'd424,  14'd1249,  14'd1406,  -14'd913,  14'd344,  -14'd213,  14'd2304,  -14'd977,  14'd863,  -14'd364,  14'd991,  14'd436,  14'd356,  

14'd1230,  -14'd96,  14'd459,  14'd505,  14'd1119,  -14'd326,  14'd739,  14'd386,  14'd635,  14'd145,  -14'd521,  -14'd201,  14'd676,  -14'd966,  14'd383,  14'd502,  
-14'd749,  -14'd328,  14'd511,  -14'd479,  -14'd997,  -14'd375,  14'd2398,  14'd784,  14'd263,  -14'd943,  14'd1023,  -14'd950,  -14'd284,  14'd569,  -14'd1524,  -14'd516,  
-14'd85,  14'd1095,  -14'd309,  14'd489,  14'd463,  -14'd17,  -14'd228,  14'd800,  14'd127,  -14'd516,  14'd101,  -14'd719,  -14'd982,  -14'd1428,  -14'd209,  -14'd554,  
14'd1209,  14'd1321,  14'd587,  14'd876,  -14'd568,  -14'd967,  -14'd559,  -14'd341,  -14'd19,  14'd324,  14'd398,  14'd799,  14'd2036,  -14'd2085,  -14'd8,  -14'd1036,  
14'd1447,  14'd1624,  -14'd1110,  14'd964,  -14'd442,  -14'd65,  -14'd114,  -14'd300,  -14'd718,  14'd1394,  -14'd888,  14'd526,  14'd816,  14'd683,  -14'd944,  14'd443,  
-14'd667,  -14'd667,  14'd639,  -14'd1248,  -14'd416,  -14'd1150,  -14'd243,  -14'd130,  14'd904,  -14'd293,  14'd1596,  -14'd229,  14'd622,  -14'd246,  14'd455,  -14'd998,  
-14'd555,  -14'd1472,  14'd350,  14'd1139,  14'd238,  -14'd780,  14'd684,  14'd897,  14'd799,  -14'd1210,  14'd704,  14'd1368,  14'd407,  14'd1364,  14'd726,  -14'd1561,  
14'd378,  -14'd1116,  14'd468,  14'd885,  -14'd976,  -14'd990,  -14'd1207,  14'd165,  14'd1116,  -14'd1177,  14'd1647,  -14'd1197,  14'd469,  -14'd176,  14'd313,  14'd285,  
-14'd1799,  14'd573,  -14'd1678,  14'd498,  14'd671,  -14'd1163,  -14'd1115,  14'd1269,  14'd494,  14'd2300,  14'd605,  14'd222,  14'd1505,  -14'd1592,  14'd818,  14'd1075,  
-14'd579,  -14'd901,  -14'd214,  14'd845,  14'd971,  14'd745,  -14'd1419,  -14'd213,  -14'd1588,  14'd3270,  14'd955,  -14'd97,  -14'd194,  -14'd937,  14'd398,  14'd894,  
-14'd449,  14'd331,  -14'd348,  14'd568,  -14'd2122,  14'd206,  14'd396,  -14'd672,  -14'd237,  -14'd725,  -14'd1499,  -14'd1547,  -14'd698,  14'd1501,  14'd19,  14'd378,  
14'd300,  -14'd304,  -14'd896,  14'd187,  -14'd753,  14'd603,  -14'd12,  14'd806,  -14'd386,  14'd68,  -14'd1237,  -14'd1510,  14'd309,  -14'd148,  14'd219,  14'd1038,  
-14'd1859,  14'd1108,  -14'd1509,  14'd357,  14'd545,  -14'd450,  14'd699,  14'd836,  14'd1794,  14'd1011,  14'd40,  -14'd686,  -14'd787,  -14'd643,  14'd1069,  14'd1240,  
-14'd2009,  14'd348,  -14'd2184,  -14'd403,  14'd1106,  -14'd50,  -14'd361,  14'd364,  -14'd216,  14'd839,  14'd1156,  14'd913,  -14'd831,  -14'd448,  -14'd68,  14'd1615,  
-14'd541,  -14'd737,  14'd1704,  -14'd52,  14'd983,  14'd1163,  14'd1331,  14'd1074,  14'd1495,  14'd768,  14'd223,  14'd1974,  -14'd205,  -14'd366,  14'd173,  -14'd454,  
14'd581,  -14'd341,  -14'd211,  14'd206,  -14'd276,  14'd547,  14'd162,  14'd819,  14'd613,  -14'd214,  -14'd1008,  -14'd666,  -14'd797,  -14'd197,  -14'd866,  14'd614,  
-14'd992,  -14'd48,  -14'd117,  -14'd272,  -14'd879,  14'd751,  14'd384,  14'd1532,  -14'd1531,  -14'd124,  14'd433,  14'd577,  -14'd139,  14'd115,  14'd889,  -14'd685,  
14'd32,  -14'd1639,  -14'd586,  -14'd189,  14'd957,  14'd265,  14'd98,  14'd708,  -14'd1093,  -14'd804,  14'd1264,  14'd1456,  14'd1155,  -14'd129,  14'd17,  14'd11,  
14'd533,  14'd1877,  -14'd447,  -14'd127,  14'd178,  14'd1903,  -14'd923,  -14'd1042,  14'd1439,  -14'd1160,  14'd391,  -14'd502,  14'd1052,  14'd629,  14'd70,  -14'd878,  
-14'd136,  -14'd189,  14'd1885,  14'd29,  -14'd312,  14'd238,  14'd598,  14'd2,  -14'd498,  -14'd898,  14'd1505,  -14'd820,  -14'd608,  14'd1047,  14'd367,  14'd100,  
14'd580,  -14'd735,  -14'd1107,  -14'd122,  -14'd509,  14'd1435,  -14'd498,  -14'd529,  -14'd270,  14'd438,  -14'd18,  14'd176,  -14'd1621,  14'd622,  14'd1020,  -14'd35,  
-14'd548,  14'd52,  -14'd760,  14'd871,  -14'd526,  14'd1770,  14'd518,  -14'd341,  14'd146,  14'd1056,  14'd180,  14'd499,  14'd131,  -14'd2052,  -14'd291,  -14'd220,  
14'd1079,  14'd341,  -14'd1587,  -14'd579,  -14'd147,  14'd565,  14'd1286,  -14'd1335,  -14'd370,  -14'd197,  14'd1772,  -14'd161,  -14'd200,  -14'd1543,  14'd458,  14'd200,  
-14'd655,  14'd804,  14'd412,  -14'd975,  14'd483,  -14'd795,  14'd1719,  -14'd340,  14'd972,  -14'd498,  -14'd196,  -14'd969,  -14'd811,  14'd1493,  14'd238,  -14'd158,  
-14'd578,  -14'd301,  -14'd855,  -14'd1243,  -14'd922,  14'd180,  -14'd531,  -14'd464,  14'd1592,  14'd119,  -14'd959,  -14'd1242,  14'd251,  14'd79,  -14'd2146,  14'd82,  

-14'd281,  -14'd574,  14'd132,  14'd427,  -14'd576,  14'd552,  14'd255,  14'd580,  -14'd681,  14'd459,  -14'd1609,  -14'd1760,  14'd334,  14'd409,  -14'd103,  14'd86,  
-14'd1705,  14'd37,  14'd614,  -14'd177,  -14'd30,  -14'd724,  -14'd305,  -14'd449,  -14'd1051,  -14'd1073,  -14'd1050,  -14'd735,  -14'd1710,  14'd1219,  14'd767,  14'd268,  
-14'd136,  -14'd427,  14'd949,  -14'd45,  -14'd726,  14'd1096,  -14'd1693,  14'd774,  14'd1398,  -14'd1082,  14'd1232,  14'd641,  14'd82,  14'd2037,  14'd355,  -14'd529,  
-14'd745,  14'd1795,  14'd1561,  -14'd725,  -14'd391,  -14'd297,  14'd664,  14'd1044,  14'd524,  -14'd285,  14'd244,  -14'd629,  -14'd98,  -14'd2247,  14'd907,  14'd1166,  
-14'd1065,  -14'd1052,  -14'd86,  14'd774,  -14'd441,  -14'd1862,  -14'd372,  -14'd835,  14'd750,  14'd211,  -14'd45,  -14'd137,  -14'd862,  14'd201,  14'd934,  -14'd1615,  
-14'd54,  14'd414,  -14'd1697,  14'd19,  14'd681,  14'd508,  -14'd1792,  -14'd1490,  -14'd501,  14'd217,  -14'd595,  -14'd221,  -14'd273,  -14'd2039,  -14'd899,  -14'd1278,  
14'd1432,  -14'd686,  14'd360,  14'd1699,  -14'd657,  -14'd396,  14'd830,  -14'd150,  -14'd1827,  14'd819,  14'd673,  -14'd52,  -14'd290,  -14'd792,  -14'd1124,  -14'd762,  
14'd350,  -14'd180,  14'd738,  -14'd1342,  -14'd1556,  -14'd106,  14'd995,  14'd195,  -14'd428,  14'd1722,  14'd264,  14'd971,  14'd618,  -14'd167,  -14'd1045,  14'd118,  
-14'd309,  -14'd499,  14'd690,  -14'd401,  -14'd1219,  -14'd249,  -14'd126,  14'd783,  -14'd1163,  14'd42,  -14'd760,  14'd148,  -14'd131,  -14'd371,  14'd765,  -14'd181,  
-14'd2222,  14'd1027,  14'd1733,  -14'd323,  -14'd991,  -14'd1817,  -14'd326,  -14'd505,  -14'd210,  14'd1190,  14'd623,  14'd264,  -14'd832,  14'd169,  14'd443,  14'd500,  
-14'd398,  14'd116,  -14'd1659,  14'd617,  -14'd163,  -14'd723,  -14'd1078,  14'd106,  14'd1928,  14'd236,  14'd2088,  14'd53,  -14'd419,  -14'd1735,  14'd258,  14'd986,  
14'd1283,  -14'd1206,  -14'd1850,  14'd687,  -14'd466,  14'd871,  -14'd445,  14'd610,  14'd731,  14'd1806,  14'd513,  14'd1388,  14'd1104,  -14'd2497,  -14'd372,  14'd858,  
14'd1805,  -14'd536,  14'd355,  14'd1183,  14'd1639,  -14'd887,  14'd823,  14'd1438,  14'd2036,  14'd1133,  14'd600,  14'd412,  14'd1789,  -14'd729,  14'd151,  14'd188,  
-14'd112,  -14'd1268,  -14'd441,  14'd883,  -14'd135,  14'd620,  -14'd95,  -14'd545,  14'd721,  14'd1333,  -14'd662,  14'd69,  -14'd930,  14'd2507,  -14'd13,  -14'd513,  
14'd3291,  14'd1311,  14'd2061,  14'd431,  -14'd2712,  14'd897,  -14'd465,  14'd390,  14'd787,  -14'd318,  -14'd772,  14'd133,  14'd1751,  -14'd1175,  14'd562,  -14'd448,  
14'd703,  -14'd1335,  14'd299,  -14'd7,  14'd2,  -14'd1059,  14'd1868,  -14'd452,  14'd3150,  14'd1344,  14'd1760,  -14'd361,  14'd386,  14'd796,  14'd491,  14'd734,  
-14'd636,  -14'd439,  -14'd495,  14'd41,  -14'd171,  14'd672,  -14'd16,  14'd661,  14'd499,  -14'd228,  14'd2648,  14'd833,  14'd1181,  14'd1092,  14'd1056,  -14'd123,  
-14'd1242,  14'd1118,  -14'd190,  14'd1699,  14'd245,  14'd1276,  14'd419,  -14'd657,  -14'd1418,  -14'd1427,  14'd1166,  14'd227,  14'd343,  -14'd117,  14'd1303,  14'd458,  
-14'd719,  14'd203,  -14'd1286,  -14'd102,  14'd614,  -14'd1143,  14'd393,  14'd33,  -14'd692,  14'd880,  -14'd1059,  -14'd2160,  14'd1294,  14'd24,  14'd292,  -14'd1183,  
14'd1720,  -14'd640,  14'd1892,  -14'd1220,  14'd1431,  -14'd1498,  -14'd1132,  14'd895,  14'd46,  14'd1212,  14'd1405,  14'd57,  14'd621,  14'd506,  -14'd1256,  -14'd277,  
14'd3,  -14'd438,  -14'd679,  -14'd17,  -14'd399,  14'd528,  14'd1042,  14'd587,  -14'd571,  -14'd616,  14'd212,  -14'd1944,  14'd1413,  14'd445,  14'd58,  14'd481,  
-14'd1874,  14'd192,  -14'd1520,  14'd60,  -14'd989,  -14'd1021,  14'd525,  -14'd1105,  -14'd307,  -14'd908,  14'd502,  -14'd1383,  14'd1008,  14'd515,  14'd252,  14'd703,  
-14'd1405,  -14'd570,  -14'd611,  -14'd628,  -14'd812,  -14'd71,  -14'd1149,  14'd200,  -14'd1825,  -14'd758,  14'd238,  -14'd1417,  -14'd1780,  14'd501,  -14'd944,  14'd1500,  
-14'd1332,  14'd337,  -14'd2335,  14'd480,  -14'd134,  -14'd128,  -14'd341,  14'd196,  14'd46,  -14'd921,  14'd526,  14'd600,  -14'd860,  -14'd1674,  14'd313,  -14'd280,  
-14'd3083,  14'd1238,  -14'd1242,  -14'd248,  -14'd697,  -14'd1935,  -14'd614,  -14'd475,  -14'd1643,  14'd158,  14'd687,  -14'd315,  -14'd1356,  14'd715,  -14'd874,  -14'd640,  

14'd189,  -14'd112,  14'd723,  -14'd103,  14'd677,  -14'd542,  -14'd755,  14'd1356,  14'd422,  14'd852,  14'd227,  14'd1826,  14'd192,  14'd1822,  14'd271,  14'd824,  
14'd329,  -14'd537,  14'd454,  14'd331,  14'd121,  14'd807,  14'd1144,  14'd492,  14'd1068,  -14'd241,  14'd1426,  14'd1365,  14'd882,  14'd1082,  -14'd39,  14'd24,  
14'd1174,  14'd395,  -14'd786,  -14'd1171,  -14'd1859,  -14'd294,  -14'd468,  14'd192,  14'd678,  14'd33,  -14'd191,  14'd102,  14'd1159,  14'd777,  -14'd1333,  -14'd1224,  
14'd970,  14'd806,  -14'd1725,  14'd618,  -14'd614,  14'd94,  14'd764,  14'd508,  -14'd1083,  14'd38,  14'd1188,  -14'd208,  14'd265,  14'd320,  -14'd644,  14'd1254,  
14'd1615,  14'd2416,  -14'd1482,  -14'd788,  14'd1283,  14'd669,  14'd512,  -14'd273,  -14'd412,  14'd622,  14'd789,  14'd128,  14'd2277,  -14'd92,  14'd129,  14'd334,  
-14'd841,  14'd1551,  14'd203,  14'd106,  14'd1105,  14'd1722,  -14'd511,  -14'd570,  14'd578,  14'd41,  -14'd671,  14'd1803,  14'd26,  14'd1288,  14'd627,  14'd571,  
14'd276,  14'd99,  14'd466,  14'd1648,  14'd397,  -14'd757,  14'd170,  -14'd509,  -14'd685,  14'd47,  14'd1473,  14'd524,  14'd224,  -14'd123,  14'd379,  -14'd711,  
-14'd1924,  -14'd1069,  14'd419,  14'd241,  -14'd710,  14'd734,  14'd786,  -14'd9,  14'd1440,  -14'd1498,  -14'd52,  -14'd946,  14'd725,  -14'd1003,  14'd233,  14'd276,  
-14'd569,  14'd476,  -14'd266,  14'd171,  14'd98,  -14'd1239,  -14'd1211,  -14'd1369,  14'd879,  14'd752,  14'd163,  14'd851,  -14'd226,  -14'd394,  -14'd404,  14'd1031,  
14'd55,  -14'd1888,  -14'd339,  14'd1148,  14'd2010,  14'd1274,  -14'd140,  14'd217,  -14'd190,  -14'd36,  -14'd950,  -14'd13,  14'd978,  -14'd2225,  -14'd959,  14'd1632,  
-14'd532,  14'd321,  14'd147,  14'd16,  14'd1465,  -14'd200,  14'd422,  -14'd976,  14'd76,  14'd588,  14'd1114,  14'd427,  14'd542,  -14'd831,  -14'd216,  14'd1375,  
-14'd227,  14'd510,  14'd886,  14'd913,  14'd560,  14'd936,  14'd912,  -14'd123,  -14'd1019,  -14'd852,  14'd574,  -14'd252,  -14'd51,  -14'd215,  14'd719,  -14'd675,  
14'd135,  -14'd1426,  14'd326,  -14'd726,  -14'd90,  14'd166,  14'd859,  -14'd1147,  14'd194,  -14'd648,  -14'd299,  14'd99,  -14'd1092,  -14'd525,  -14'd632,  -14'd596,  
-14'd1162,  -14'd1192,  -14'd1930,  14'd399,  -14'd112,  -14'd448,  14'd82,  -14'd1042,  14'd798,  -14'd377,  -14'd276,  14'd72,  14'd155,  -14'd117,  14'd960,  -14'd61,  
-14'd739,  -14'd790,  -14'd812,  -14'd83,  14'd541,  14'd257,  -14'd75,  14'd77,  -14'd900,  14'd1474,  14'd1647,  14'd186,  14'd571,  14'd1272,  14'd1296,  14'd1307,  
14'd75,  14'd658,  14'd42,  -14'd1482,  -14'd1460,  -14'd304,  14'd883,  -14'd1026,  -14'd727,  14'd301,  -14'd890,  14'd239,  -14'd348,  -14'd581,  -14'd523,  14'd1091,  
14'd1991,  14'd169,  14'd79,  14'd618,  14'd1238,  -14'd1198,  14'd211,  -14'd902,  -14'd1632,  14'd93,  -14'd1560,  14'd348,  14'd592,  14'd929,  14'd750,  -14'd123,  
14'd326,  14'd1596,  14'd819,  -14'd201,  14'd1022,  -14'd54,  14'd905,  -14'd776,  14'd1112,  -14'd381,  14'd1482,  -14'd1421,  -14'd602,  -14'd1361,  14'd390,  -14'd32,  
14'd107,  -14'd251,  -14'd1234,  14'd1457,  -14'd292,  14'd185,  14'd211,  -14'd1606,  -14'd408,  14'd1479,  -14'd533,  -14'd545,  -14'd187,  -14'd1272,  14'd678,  14'd123,  
-14'd1665,  -14'd281,  14'd1277,  14'd976,  14'd325,  -14'd918,  -14'd73,  14'd477,  -14'd735,  14'd731,  -14'd344,  14'd1561,  -14'd635,  14'd974,  -14'd1283,  14'd127,  
14'd721,  -14'd151,  -14'd1249,  -14'd161,  -14'd742,  -14'd585,  -14'd1768,  -14'd1061,  -14'd1245,  14'd1287,  -14'd268,  14'd53,  14'd82,  14'd2580,  -14'd1047,  -14'd399,  
14'd31,  14'd836,  -14'd842,  14'd256,  -14'd435,  -14'd391,  -14'd1993,  -14'd27,  14'd467,  -14'd643,  -14'd1090,  -14'd751,  14'd59,  14'd369,  14'd344,  -14'd575,  
14'd954,  -14'd152,  -14'd2013,  -14'd528,  -14'd554,  14'd915,  -14'd50,  14'd1057,  -14'd555,  -14'd1805,  14'd1043,  -14'd502,  -14'd606,  -14'd705,  14'd745,  14'd635,  
14'd1071,  14'd677,  -14'd511,  14'd635,  -14'd616,  14'd121,  -14'd580,  14'd775,  14'd64,  -14'd1595,  14'd142,  14'd429,  14'd433,  -14'd55,  -14'd227,  14'd254,  
-14'd1281,  -14'd631,  -14'd1586,  -14'd468,  -14'd435,  -14'd543,  14'd248,  14'd268,  -14'd1567,  -14'd3343,  -14'd669,  -14'd1706,  -14'd1303,  -14'd159,  -14'd152,  -14'd894,  

14'd888,  14'd809,  14'd1799,  14'd1259,  14'd849,  14'd315,  14'd1102,  14'd551,  14'd1263,  14'd908,  14'd579,  -14'd694,  14'd647,  14'd1918,  14'd1091,  -14'd1551,  
-14'd1455,  -14'd1480,  14'd1064,  14'd1078,  14'd976,  -14'd6,  -14'd621,  -14'd670,  -14'd509,  14'd1194,  14'd250,  14'd324,  -14'd127,  -14'd160,  -14'd129,  14'd175,  
-14'd614,  -14'd65,  -14'd107,  14'd299,  -14'd703,  14'd627,  14'd277,  14'd592,  14'd48,  14'd189,  14'd1095,  14'd1604,  14'd207,  -14'd2521,  -14'd482,  -14'd1664,  
14'd798,  -14'd99,  -14'd144,  -14'd288,  14'd1635,  -14'd1255,  -14'd1308,  14'd155,  -14'd886,  14'd1141,  -14'd66,  -14'd920,  14'd1245,  -14'd2705,  -14'd1685,  14'd1178,  
14'd1535,  -14'd1745,  -14'd1538,  -14'd49,  -14'd993,  14'd118,  -14'd1094,  14'd1505,  -14'd350,  14'd362,  -14'd513,  -14'd1648,  -14'd253,  -14'd933,  -14'd365,  -14'd476,  
-14'd711,  14'd1131,  -14'd1166,  14'd1136,  14'd915,  14'd406,  -14'd1013,  14'd1255,  14'd564,  14'd599,  14'd1289,  14'd271,  -14'd306,  -14'd100,  14'd1744,  -14'd358,  
-14'd375,  -14'd463,  14'd530,  14'd738,  14'd607,  14'd558,  14'd179,  14'd651,  14'd507,  14'd852,  14'd403,  14'd792,  -14'd687,  -14'd1150,  -14'd529,  -14'd868,  
-14'd2658,  14'd969,  -14'd1550,  -14'd582,  14'd1251,  -14'd1526,  14'd1051,  14'd1201,  -14'd126,  14'd42,  14'd538,  14'd318,  14'd237,  -14'd310,  14'd388,  -14'd170,  
14'd610,  14'd45,  -14'd21,  14'd727,  14'd370,  -14'd85,  -14'd1525,  -14'd184,  -14'd993,  14'd300,  14'd8,  -14'd12,  14'd605,  -14'd12,  14'd419,  -14'd81,  
14'd1906,  -14'd448,  -14'd1835,  -14'd34,  -14'd742,  14'd12,  -14'd861,  14'd37,  14'd91,  14'd1452,  14'd654,  14'd423,  14'd1093,  -14'd1963,  14'd525,  14'd1094,  
14'd646,  14'd170,  -14'd354,  14'd383,  14'd1704,  -14'd697,  -14'd446,  14'd168,  -14'd738,  -14'd1688,  14'd822,  14'd360,  14'd205,  -14'd36,  -14'd245,  -14'd434,  
-14'd18,  14'd120,  -14'd231,  -14'd968,  -14'd1016,  -14'd544,  -14'd918,  -14'd1477,  -14'd275,  -14'd31,  14'd1611,  -14'd206,  14'd74,  -14'd1540,  14'd1075,  14'd396,  
14'd137,  -14'd731,  14'd555,  14'd480,  -14'd985,  -14'd491,  -14'd465,  14'd621,  -14'd153,  -14'd1036,  14'd2736,  -14'd1031,  -14'd506,  14'd1311,  14'd1435,  14'd488,  
-14'd127,  14'd842,  14'd212,  14'd1092,  14'd229,  14'd53,  14'd270,  -14'd4,  14'd1152,  -14'd1298,  14'd264,  14'd425,  14'd1245,  -14'd452,  -14'd285,  14'd764,  
-14'd2454,  -14'd901,  14'd713,  14'd1791,  14'd504,  14'd673,  14'd27,  -14'd431,  14'd419,  14'd521,  14'd876,  14'd261,  14'd1527,  14'd231,  14'd1417,  -14'd332,  
14'd773,  14'd537,  14'd313,  -14'd566,  14'd418,  -14'd957,  14'd241,  14'd462,  -14'd1083,  -14'd115,  14'd1226,  14'd58,  14'd762,  -14'd518,  14'd59,  -14'd267,  
-14'd793,  14'd142,  -14'd1705,  -14'd1256,  -14'd209,  -14'd1941,  -14'd166,  -14'd584,  -14'd331,  -14'd304,  14'd532,  14'd247,  14'd270,  14'd207,  -14'd1816,  14'd722,  
14'd1157,  14'd1498,  14'd15,  -14'd1645,  14'd267,  -14'd1358,  14'd335,  -14'd101,  14'd390,  14'd835,  -14'd44,  -14'd576,  -14'd414,  14'd1279,  -14'd124,  -14'd91,  
14'd1382,  14'd1814,  14'd1646,  -14'd1157,  -14'd11,  -14'd266,  14'd286,  14'd1203,  14'd1505,  14'd554,  14'd640,  14'd1211,  -14'd1240,  -14'd105,  14'd1473,  -14'd821,  
14'd277,  14'd710,  -14'd115,  14'd1053,  14'd1377,  14'd456,  -14'd172,  14'd234,  14'd516,  -14'd121,  14'd1341,  -14'd1455,  14'd139,  14'd735,  -14'd537,  14'd1243,  
-14'd43,  14'd170,  -14'd422,  -14'd1763,  14'd48,  -14'd547,  14'd867,  -14'd1637,  14'd326,  -14'd2087,  -14'd1375,  14'd586,  -14'd2061,  -14'd1587,  14'd207,  14'd683,  
-14'd560,  -14'd343,  -14'd1800,  -14'd134,  -14'd52,  -14'd207,  14'd1273,  -14'd789,  14'd1596,  -14'd770,  -14'd1013,  14'd527,  -14'd703,  14'd303,  -14'd411,  14'd63,  
14'd1019,  -14'd633,  14'd1220,  -14'd486,  14'd757,  -14'd211,  14'd1355,  -14'd1268,  14'd3097,  14'd366,  -14'd193,  -14'd105,  -14'd893,  14'd1052,  -14'd462,  -14'd1123,  
-14'd593,  14'd347,  14'd633,  -14'd709,  -14'd21,  -14'd644,  -14'd812,  14'd862,  14'd27,  14'd33,  -14'd944,  -14'd786,  -14'd64,  14'd1336,  14'd149,  -14'd555,  
-14'd842,  14'd236,  14'd427,  14'd466,  -14'd953,  14'd234,  -14'd841,  -14'd83,  14'd397,  14'd1894,  14'd264,  -14'd333,  -14'd1231,  -14'd422,  -14'd1466,  -14'd351,  

14'd396,  14'd1836,  14'd502,  -14'd417,  -14'd725,  14'd105,  14'd2322,  -14'd567,  14'd107,  -14'd117,  -14'd136,  14'd2129,  -14'd1721,  14'd1595,  -14'd1628,  14'd325,  
14'd20,  14'd760,  -14'd796,  -14'd448,  -14'd1656,  -14'd625,  14'd1988,  14'd225,  14'd1099,  -14'd330,  -14'd196,  14'd170,  -14'd1231,  14'd4,  14'd353,  14'd275,  
14'd1723,  14'd610,  -14'd29,  -14'd1158,  14'd837,  -14'd997,  -14'd388,  14'd614,  14'd1063,  -14'd12,  14'd78,  14'd54,  14'd389,  14'd93,  14'd46,  -14'd520,  
-14'd74,  -14'd228,  14'd89,  14'd336,  -14'd109,  14'd1358,  14'd522,  14'd44,  14'd533,  14'd537,  -14'd400,  -14'd687,  14'd976,  -14'd739,  -14'd256,  -14'd5,  
-14'd2154,  14'd1505,  14'd790,  -14'd283,  -14'd1076,  14'd1079,  -14'd518,  14'd54,  14'd438,  -14'd308,  14'd1451,  14'd72,  14'd1062,  14'd1552,  14'd1236,  14'd1370,  
-14'd1161,  -14'd1437,  14'd262,  -14'd1104,  -14'd803,  -14'd419,  14'd1163,  14'd320,  14'd1021,  -14'd486,  -14'd142,  -14'd392,  -14'd1407,  14'd375,  14'd519,  14'd307,  
14'd892,  -14'd338,  14'd430,  -14'd1548,  14'd407,  14'd128,  -14'd1164,  -14'd619,  14'd916,  14'd445,  -14'd636,  -14'd452,  -14'd374,  14'd1182,  14'd794,  14'd65,  
-14'd1148,  -14'd877,  -14'd39,  -14'd862,  14'd457,  -14'd535,  14'd240,  14'd1052,  -14'd624,  14'd704,  14'd1077,  14'd581,  -14'd1707,  -14'd555,  14'd174,  -14'd801,  
-14'd281,  -14'd59,  -14'd68,  -14'd537,  14'd899,  14'd189,  -14'd300,  -14'd637,  -14'd876,  14'd2272,  -14'd380,  -14'd57,  14'd89,  -14'd1009,  14'd134,  -14'd238,  
-14'd1285,  -14'd1148,  -14'd326,  -14'd326,  -14'd1082,  -14'd1451,  14'd813,  14'd287,  14'd119,  14'd503,  -14'd605,  -14'd427,  -14'd641,  -14'd559,  -14'd1714,  14'd830,  
-14'd658,  14'd980,  -14'd292,  -14'd90,  14'd314,  14'd1364,  -14'd722,  14'd296,  -14'd1518,  14'd1642,  -14'd1045,  -14'd277,  14'd140,  -14'd68,  14'd396,  14'd217,  
14'd1895,  14'd752,  14'd285,  14'd157,  -14'd95,  14'd429,  -14'd5,  14'd981,  -14'd139,  -14'd326,  14'd534,  -14'd851,  -14'd1899,  14'd1670,  14'd257,  -14'd1443,  
-14'd426,  14'd944,  -14'd863,  -14'd76,  14'd1546,  14'd572,  14'd341,  14'd601,  14'd1505,  -14'd722,  -14'd395,  14'd1364,  -14'd796,  -14'd909,  -14'd678,  -14'd1155,  
14'd289,  14'd272,  -14'd1117,  -14'd2435,  14'd899,  14'd778,  14'd461,  -14'd1116,  14'd1659,  14'd1085,  -14'd407,  -14'd1072,  14'd123,  -14'd108,  -14'd259,  -14'd295,  
-14'd1329,  -14'd823,  -14'd785,  14'd1191,  -14'd1670,  14'd1054,  -14'd1022,  -14'd314,  14'd803,  14'd1087,  14'd388,  -14'd105,  -14'd1741,  -14'd156,  -14'd150,  14'd1542,  
14'd211,  -14'd195,  14'd1497,  14'd765,  -14'd157,  14'd308,  -14'd137,  -14'd275,  -14'd732,  -14'd312,  -14'd1770,  14'd1110,  -14'd576,  14'd489,  -14'd25,  14'd725,  
14'd1186,  14'd357,  -14'd767,  14'd1310,  -14'd268,  14'd418,  -14'd799,  14'd216,  14'd1885,  -14'd707,  -14'd1206,  14'd703,  14'd885,  14'd610,  14'd1574,  14'd577,  
-14'd664,  -14'd635,  -14'd76,  14'd127,  -14'd183,  14'd354,  14'd1327,  14'd1562,  -14'd1155,  -14'd1187,  14'd17,  -14'd309,  -14'd1894,  14'd776,  14'd925,  -14'd252,  
-14'd77,  14'd610,  -14'd545,  14'd159,  14'd844,  14'd622,  -14'd298,  -14'd1452,  -14'd540,  -14'd215,  -14'd855,  14'd1094,  -14'd58,  14'd1996,  14'd85,  -14'd748,  
-14'd716,  14'd538,  14'd1288,  14'd507,  -14'd408,  14'd642,  14'd1167,  -14'd953,  14'd1284,  14'd193,  -14'd414,  -14'd45,  -14'd1029,  14'd971,  -14'd412,  -14'd154,  
-14'd1627,  -14'd1126,  -14'd608,  14'd986,  14'd741,  14'd2018,  -14'd727,  14'd1948,  14'd596,  14'd295,  -14'd788,  -14'd874,  14'd1021,  -14'd1152,  14'd65,  14'd655,  
14'd57,  14'd1175,  14'd173,  14'd747,  14'd2268,  -14'd14,  -14'd1015,  14'd2067,  -14'd667,  -14'd1095,  14'd1793,  -14'd903,  -14'd26,  -14'd822,  14'd1358,  -14'd36,  
-14'd691,  -14'd700,  -14'd837,  14'd1221,  14'd127,  14'd1236,  -14'd394,  14'd1339,  14'd444,  14'd1121,  14'd1069,  14'd194,  14'd996,  -14'd209,  14'd74,  14'd504,  
14'd86,  14'd1425,  -14'd1095,  14'd1660,  -14'd416,  14'd1590,  14'd4,  14'd705,  14'd258,  14'd1143,  -14'd1062,  14'd2096,  14'd1354,  -14'd121,  14'd129,  -14'd520,  
14'd1955,  14'd442,  14'd655,  14'd1516,  14'd599,  14'd291,  14'd515,  14'd1724,  14'd2783,  14'd432,  14'd722,  14'd1399,  -14'd51,  14'd973,  -14'd310,  -14'd321,  

-14'd316,  -14'd168,  14'd346,  14'd145,  -14'd167,  14'd465,  14'd1413,  14'd985,  -14'd1259,  -14'd767,  -14'd245,  -14'd123,  -14'd375,  -14'd1153,  14'd166,  -14'd320,  
14'd198,  -14'd1276,  14'd133,  -14'd1107,  14'd345,  -14'd216,  -14'd1035,  -14'd1730,  -14'd1630,  -14'd842,  -14'd505,  -14'd1122,  14'd151,  14'd243,  -14'd1607,  -14'd1231,  
-14'd65,  14'd237,  14'd465,  14'd750,  -14'd1195,  -14'd419,  -14'd726,  -14'd235,  -14'd78,  14'd178,  -14'd130,  -14'd1920,  14'd83,  14'd675,  -14'd1091,  14'd843,  
-14'd1276,  -14'd609,  -14'd1245,  14'd275,  14'd488,  -14'd1545,  -14'd172,  -14'd589,  14'd298,  -14'd754,  -14'd349,  14'd175,  -14'd187,  14'd58,  -14'd265,  -14'd123,  
-14'd87,  14'd241,  -14'd937,  -14'd809,  14'd17,  -14'd292,  -14'd292,  14'd132,  14'd267,  14'd975,  -14'd686,  14'd130,  14'd246,  -14'd662,  -14'd1032,  -14'd1032,  
-14'd650,  -14'd590,  -14'd374,  -14'd649,  -14'd1536,  14'd1048,  -14'd996,  14'd901,  14'd915,  -14'd43,  -14'd730,  -14'd1094,  14'd993,  -14'd473,  14'd799,  -14'd1162,  
-14'd64,  14'd107,  14'd42,  14'd893,  14'd675,  14'd1041,  -14'd1086,  -14'd1814,  -14'd275,  14'd1094,  14'd967,  -14'd454,  14'd603,  14'd600,  14'd604,  -14'd1215,  
14'd1121,  14'd702,  -14'd665,  -14'd1371,  14'd380,  14'd602,  -14'd190,  14'd248,  -14'd437,  -14'd81,  -14'd1045,  14'd406,  14'd419,  14'd589,  -14'd795,  -14'd1063,  
-14'd540,  -14'd190,  -14'd1029,  14'd2,  14'd130,  -14'd905,  -14'd1195,  -14'd1079,  -14'd396,  14'd284,  -14'd987,  -14'd341,  -14'd1089,  -14'd326,  14'd371,  -14'd506,  
14'd1091,  14'd452,  14'd1374,  -14'd838,  -14'd739,  14'd646,  -14'd459,  -14'd443,  -14'd808,  14'd552,  -14'd471,  -14'd1323,  -14'd1218,  14'd603,  -14'd1015,  14'd342,  
-14'd755,  -14'd1070,  -14'd1177,  14'd239,  -14'd634,  14'd431,  -14'd617,  -14'd1631,  14'd776,  -14'd793,  -14'd1647,  -14'd266,  -14'd337,  -14'd282,  -14'd281,  -14'd840,  
14'd353,  -14'd775,  -14'd62,  -14'd390,  -14'd1307,  -14'd298,  14'd364,  -14'd750,  -14'd762,  14'd677,  -14'd591,  -14'd975,  -14'd997,  -14'd616,  14'd484,  -14'd843,  
14'd429,  -14'd220,  -14'd1419,  14'd455,  -14'd554,  -14'd1585,  -14'd38,  14'd510,  -14'd306,  -14'd730,  14'd245,  -14'd1700,  -14'd639,  -14'd389,  14'd826,  -14'd56,  
14'd352,  -14'd1090,  -14'd1463,  14'd1222,  -14'd696,  -14'd141,  -14'd152,  -14'd637,  -14'd1579,  14'd19,  -14'd907,  -14'd1233,  -14'd530,  -14'd247,  14'd888,  -14'd240,  
14'd505,  14'd335,  -14'd961,  14'd336,  -14'd23,  -14'd362,  -14'd770,  -14'd132,  -14'd920,  14'd828,  -14'd450,  -14'd381,  14'd213,  14'd1376,  -14'd550,  14'd1020,  
-14'd13,  14'd419,  -14'd886,  -14'd693,  -14'd258,  -14'd343,  14'd253,  -14'd393,  14'd466,  -14'd996,  14'd744,  -14'd523,  -14'd841,  14'd6,  -14'd452,  -14'd192,  
14'd867,  -14'd908,  14'd490,  -14'd33,  -14'd1250,  -14'd1105,  -14'd265,  14'd155,  -14'd48,  -14'd1585,  -14'd536,  14'd407,  -14'd29,  -14'd483,  -14'd1852,  -14'd577,  
14'd928,  -14'd509,  -14'd1128,  -14'd820,  14'd579,  -14'd717,  -14'd581,  -14'd541,  14'd263,  -14'd1646,  -14'd860,  -14'd282,  14'd521,  -14'd1720,  14'd679,  14'd335,  
14'd40,  -14'd591,  14'd337,  -14'd382,  -14'd105,  14'd975,  14'd576,  -14'd933,  -14'd783,  14'd360,  -14'd498,  14'd67,  14'd161,  -14'd485,  -14'd1387,  -14'd777,  
14'd105,  -14'd404,  -14'd822,  -14'd1675,  14'd468,  14'd491,  -14'd1671,  -14'd1749,  -14'd86,  14'd712,  -14'd167,  14'd693,  -14'd1361,  -14'd46,  14'd22,  14'd196,  
-14'd561,  -14'd913,  -14'd1797,  -14'd461,  -14'd1442,  -14'd1553,  -14'd301,  -14'd1492,  -14'd1163,  -14'd851,  -14'd172,  -14'd338,  -14'd587,  14'd802,  -14'd638,  -14'd209,  
-14'd964,  14'd148,  -14'd286,  -14'd1636,  -14'd1168,  -14'd1164,  14'd212,  -14'd1236,  14'd577,  -14'd591,  -14'd947,  14'd253,  -14'd875,  -14'd534,  -14'd1669,  14'd30,  
14'd1017,  -14'd342,  -14'd234,  14'd374,  -14'd75,  -14'd169,  -14'd717,  14'd164,  14'd688,  14'd38,  -14'd447,  -14'd1430,  -14'd113,  -14'd1059,  14'd61,  -14'd73,  
14'd1305,  14'd505,  14'd811,  -14'd1540,  -14'd336,  14'd146,  -14'd1071,  -14'd557,  -14'd1218,  14'd656,  -14'd1542,  14'd211,  -14'd1496,  14'd631,  -14'd1277,  -14'd492,  
14'd1364,  14'd1049,  -14'd169,  -14'd957,  -14'd360,  -14'd1010,  14'd328,  -14'd45,  14'd470,  -14'd45,  14'd1222,  -14'd1092,  -14'd342,  14'd91,  -14'd31,  -14'd1047,  

14'd591,  -14'd1368,  14'd736,  -14'd598,  -14'd1053,  -14'd205,  -14'd836,  -14'd657,  -14'd124,  14'd1767,  -14'd1479,  -14'd1516,  -14'd1542,  -14'd645,  -14'd1954,  -14'd403,  
-14'd1040,  -14'd2286,  -14'd618,  -14'd51,  -14'd274,  14'd1230,  14'd131,  -14'd6,  -14'd2222,  -14'd2,  -14'd1249,  -14'd1846,  -14'd1185,  -14'd2229,  -14'd1080,  14'd226,  
-14'd438,  14'd601,  -14'd51,  14'd669,  -14'd1384,  14'd492,  -14'd2365,  -14'd528,  -14'd408,  -14'd913,  -14'd2072,  14'd562,  -14'd482,  14'd270,  -14'd1768,  -14'd788,  
-14'd276,  14'd782,  -14'd40,  14'd122,  14'd229,  14'd1892,  -14'd492,  -14'd1245,  14'd665,  -14'd427,  -14'd1239,  -14'd1182,  -14'd996,  -14'd1498,  -14'd326,  14'd436,  
14'd1774,  14'd1295,  14'd702,  14'd1344,  -14'd1095,  14'd764,  -14'd508,  14'd755,  14'd863,  -14'd654,  -14'd257,  -14'd1308,  -14'd619,  -14'd555,  14'd224,  14'd466,  
-14'd1476,  -14'd961,  -14'd2104,  14'd210,  -14'd570,  -14'd1033,  -14'd2186,  -14'd1462,  -14'd418,  14'd708,  14'd1834,  14'd1488,  14'd209,  -14'd273,  -14'd270,  -14'd1207,  
-14'd550,  -14'd712,  14'd195,  14'd846,  14'd176,  14'd746,  -14'd614,  -14'd1014,  14'd874,  14'd745,  14'd1925,  -14'd1064,  14'd736,  -14'd189,  -14'd114,  -14'd0,  
14'd1012,  14'd430,  14'd396,  14'd1045,  14'd150,  14'd528,  -14'd110,  14'd1770,  14'd232,  14'd869,  -14'd11,  -14'd162,  14'd1634,  14'd1381,  14'd336,  -14'd215,  
14'd2035,  14'd23,  -14'd186,  -14'd268,  14'd538,  14'd1420,  -14'd663,  14'd282,  14'd1606,  -14'd209,  14'd2541,  -14'd599,  14'd742,  14'd984,  -14'd255,  -14'd4,  
14'd456,  14'd537,  14'd596,  -14'd273,  14'd1643,  -14'd1364,  -14'd1413,  -14'd110,  -14'd536,  14'd2171,  -14'd1575,  14'd1024,  -14'd613,  14'd1855,  14'd1,  14'd482,  
-14'd1362,  14'd221,  -14'd1758,  14'd158,  -14'd495,  14'd886,  14'd1447,  14'd504,  14'd2397,  -14'd379,  14'd1687,  -14'd1195,  -14'd82,  14'd701,  14'd1425,  14'd1218,  
-14'd672,  14'd85,  -14'd546,  14'd340,  -14'd110,  -14'd601,  14'd408,  -14'd1228,  14'd1441,  -14'd101,  14'd972,  -14'd949,  -14'd1840,  14'd1925,  14'd1659,  14'd1092,  
-14'd423,  -14'd754,  -14'd700,  -14'd1038,  14'd112,  -14'd1908,  -14'd857,  14'd550,  -14'd1832,  -14'd420,  -14'd645,  -14'd1851,  -14'd220,  14'd461,  14'd1485,  14'd1146,  
14'd435,  14'd649,  -14'd1060,  -14'd430,  -14'd771,  -14'd1178,  -14'd2105,  -14'd324,  -14'd1037,  -14'd372,  14'd40,  -14'd842,  -14'd1928,  14'd1336,  14'd358,  14'd276,  
14'd1047,  -14'd335,  14'd1606,  -14'd705,  -14'd789,  -14'd1154,  14'd148,  -14'd1626,  14'd588,  14'd1862,  -14'd1636,  14'd1649,  -14'd1277,  14'd397,  14'd389,  14'd675,  
-14'd269,  -14'd1869,  14'd1236,  -14'd151,  -14'd610,  -14'd756,  14'd203,  -14'd466,  -14'd1290,  14'd156,  14'd1786,  -14'd1376,  -14'd1419,  -14'd1410,  -14'd1360,  -14'd116,  
14'd487,  -14'd721,  -14'd870,  14'd627,  -14'd1015,  -14'd1411,  -14'd569,  14'd211,  -14'd1684,  -14'd1547,  14'd359,  -14'd1677,  -14'd80,  -14'd312,  -14'd1032,  14'd255,  
14'd189,  14'd1554,  -14'd461,  -14'd108,  -14'd1140,  -14'd659,  14'd798,  14'd554,  14'd2022,  14'd1002,  -14'd1081,  -14'd953,  -14'd1690,  -14'd621,  -14'd770,  -14'd1225,  
14'd457,  14'd954,  14'd205,  -14'd842,  -14'd1762,  14'd278,  14'd96,  14'd585,  14'd587,  14'd54,  14'd123,  14'd704,  -14'd894,  14'd508,  -14'd288,  -14'd982,  
14'd1557,  -14'd471,  14'd476,  -14'd243,  -14'd1335,  14'd1207,  14'd443,  14'd1022,  14'd805,  -14'd180,  14'd905,  14'd160,  14'd1253,  14'd851,  14'd1289,  14'd464,  
-14'd1563,  14'd1713,  -14'd1984,  -14'd1528,  14'd1129,  -14'd1217,  -14'd1832,  -14'd1565,  -14'd613,  -14'd1487,  -14'd921,  14'd655,  -14'd325,  14'd730,  -14'd640,  -14'd304,  
-14'd341,  14'd687,  14'd341,  -14'd2425,  -14'd317,  -14'd1108,  -14'd856,  -14'd1495,  -14'd1421,  -14'd662,  14'd349,  -14'd221,  -14'd1169,  14'd318,  -14'd28,  -14'd1296,  
14'd1168,  -14'd797,  14'd1360,  -14'd115,  -14'd1156,  -14'd730,  -14'd966,  -14'd215,  14'd1374,  -14'd228,  -14'd2273,  -14'd28,  -14'd1898,  14'd125,  14'd556,  -14'd1351,  
14'd1885,  -14'd1774,  14'd1040,  14'd27,  14'd1063,  14'd314,  -14'd602,  -14'd1021,  14'd78,  14'd1422,  14'd585,  -14'd24,  14'd317,  14'd229,  14'd299,  -14'd37,  
14'd1168,  -14'd682,  -14'd1485,  -14'd278,  14'd272,  14'd1123,  -14'd61,  14'd1033,  14'd687,  -14'd5,  14'd622,  14'd629,  -14'd68,  -14'd700,  14'd2122,  14'd1077,  

-14'd267,  -14'd1175,  -14'd526,  14'd1844,  14'd364,  14'd1332,  14'd617,  14'd1177,  14'd935,  14'd688,  14'd1633,  -14'd28,  14'd852,  -14'd577,  14'd588,  -14'd18,  
-14'd1614,  -14'd809,  14'd1381,  14'd1710,  14'd163,  14'd833,  -14'd657,  14'd1089,  14'd416,  14'd1922,  14'd1397,  -14'd1230,  14'd1146,  -14'd483,  14'd1958,  -14'd747,  
-14'd829,  -14'd1817,  -14'd410,  -14'd5,  -14'd1271,  14'd250,  -14'd872,  14'd970,  -14'd126,  14'd242,  -14'd217,  14'd340,  14'd1391,  -14'd2986,  -14'd434,  -14'd307,  
14'd768,  14'd364,  -14'd176,  14'd676,  14'd606,  14'd553,  -14'd756,  -14'd549,  -14'd635,  14'd107,  -14'd911,  14'd757,  14'd1511,  -14'd3021,  -14'd607,  -14'd204,  
-14'd70,  14'd314,  14'd180,  14'd262,  -14'd555,  14'd409,  -14'd509,  -14'd246,  -14'd943,  -14'd932,  -14'd1163,  -14'd330,  14'd1879,  -14'd307,  -14'd111,  14'd582,  
-14'd654,  -14'd852,  -14'd660,  14'd550,  -14'd389,  -14'd560,  -14'd2066,  14'd258,  -14'd416,  -14'd524,  14'd988,  14'd13,  14'd120,  14'd1385,  14'd360,  -14'd193,  
-14'd297,  14'd340,  -14'd372,  14'd493,  14'd25,  14'd196,  -14'd170,  -14'd213,  14'd899,  -14'd1346,  14'd363,  14'd501,  14'd680,  14'd755,  -14'd228,  -14'd534,  
-14'd1941,  14'd886,  -14'd391,  14'd352,  -14'd932,  14'd690,  -14'd1562,  -14'd569,  14'd2818,  14'd183,  14'd713,  14'd171,  14'd149,  -14'd1229,  -14'd305,  14'd715,  
-14'd126,  -14'd532,  -14'd1378,  -14'd286,  -14'd947,  -14'd837,  -14'd1663,  14'd844,  14'd851,  14'd1617,  -14'd558,  14'd579,  14'd1747,  -14'd2326,  -14'd613,  14'd1038,  
14'd516,  14'd202,  -14'd1001,  -14'd201,  14'd1566,  14'd261,  14'd505,  14'd515,  14'd889,  14'd601,  14'd1094,  -14'd598,  14'd203,  -14'd388,  -14'd1489,  14'd528,  
-14'd474,  -14'd40,  14'd1212,  14'd349,  -14'd685,  14'd603,  -14'd165,  14'd819,  14'd2,  -14'd178,  -14'd319,  -14'd1294,  14'd413,  14'd418,  -14'd1364,  14'd388,  
14'd356,  14'd13,  14'd1525,  -14'd519,  -14'd320,  -14'd788,  14'd1146,  14'd482,  -14'd683,  -14'd1371,  14'd941,  -14'd841,  -14'd595,  -14'd640,  14'd786,  14'd472,  
14'd651,  14'd313,  14'd565,  -14'd747,  -14'd1031,  -14'd375,  14'd554,  -14'd366,  -14'd739,  14'd201,  -14'd154,  -14'd1252,  -14'd36,  14'd73,  -14'd232,  14'd1741,  
-14'd1058,  14'd1249,  -14'd184,  14'd261,  14'd176,  14'd1290,  -14'd153,  14'd827,  14'd1047,  14'd72,  -14'd354,  -14'd479,  14'd483,  -14'd135,  14'd496,  14'd1001,  
-14'd3148,  -14'd393,  -14'd1022,  -14'd332,  -14'd112,  -14'd1798,  14'd363,  14'd101,  14'd238,  -14'd226,  14'd1659,  14'd789,  -14'd1064,  -14'd446,  14'd1545,  14'd467,  
14'd277,  -14'd139,  14'd29,  -14'd298,  -14'd1155,  -14'd625,  14'd1143,  -14'd1705,  14'd907,  -14'd47,  14'd430,  -14'd393,  -14'd226,  14'd187,  -14'd1470,  -14'd1540,  
-14'd630,  -14'd561,  -14'd722,  -14'd975,  -14'd468,  14'd264,  -14'd565,  14'd839,  -14'd1359,  14'd2043,  14'd1425,  14'd648,  -14'd508,  14'd3,  -14'd5,  14'd187,  
-14'd105,  14'd376,  -14'd724,  14'd679,  14'd281,  14'd8,  -14'd1203,  14'd928,  14'd876,  -14'd1000,  -14'd801,  -14'd425,  14'd267,  14'd1107,  -14'd16,  -14'd1450,  
14'd300,  -14'd165,  14'd1230,  -14'd208,  14'd431,  14'd368,  -14'd2,  -14'd359,  -14'd1018,  -14'd821,  14'd930,  14'd51,  -14'd1099,  -14'd226,  -14'd1062,  -14'd767,  
14'd653,  14'd1203,  14'd966,  -14'd727,  -14'd80,  -14'd281,  14'd754,  14'd1089,  14'd189,  -14'd34,  14'd480,  -14'd41,  -14'd437,  14'd1218,  -14'd227,  -14'd1347,  
14'd588,  -14'd321,  -14'd204,  14'd1299,  -14'd1133,  -14'd1254,  14'd1843,  14'd61,  14'd1925,  14'd540,  14'd531,  14'd190,  -14'd649,  -14'd2006,  14'd58,  14'd1052,  
-14'd497,  14'd29,  -14'd1453,  14'd1125,  -14'd423,  14'd330,  14'd889,  -14'd290,  14'd423,  -14'd665,  14'd28,  -14'd299,  -14'd640,  14'd462,  -14'd1208,  14'd923,  
14'd704,  -14'd327,  14'd1159,  -14'd1168,  -14'd171,  -14'd785,  -14'd214,  14'd448,  14'd2227,  -14'd208,  14'd702,  14'd180,  -14'd324,  14'd218,  -14'd1480,  -14'd872,  
14'd468,  14'd1361,  14'd229,  14'd571,  -14'd660,  -14'd348,  -14'd95,  -14'd144,  14'd1779,  -14'd141,  14'd625,  -14'd1087,  14'd519,  14'd407,  -14'd94,  -14'd204,  
14'd286,  14'd635,  -14'd202,  -14'd1844,  -14'd1193,  -14'd1049,  -14'd261,  -14'd123,  -14'd63,  -14'd950,  -14'd935,  -14'd1003,  -14'd427,  14'd828,  -14'd409,  -14'd480,  

-14'd1385,  14'd476,  14'd1202,  14'd1623,  14'd107,  14'd526,  -14'd2384,  14'd2371,  -14'd494,  14'd2213,  -14'd1996,  14'd241,  14'd969,  -14'd821,  -14'd241,  -14'd83,  
-14'd57,  14'd952,  14'd3490,  14'd557,  14'd1315,  -14'd135,  -14'd182,  14'd1080,  14'd1121,  -14'd51,  -14'd843,  -14'd387,  -14'd354,  14'd1934,  -14'd552,  -14'd1544,  
14'd695,  14'd291,  14'd2966,  14'd694,  -14'd1402,  14'd402,  14'd1045,  -14'd612,  14'd232,  -14'd984,  -14'd205,  -14'd288,  -14'd611,  14'd2043,  14'd801,  -14'd1311,  
14'd208,  -14'd9,  14'd285,  14'd1231,  -14'd317,  -14'd1030,  14'd509,  14'd478,  -14'd830,  -14'd19,  14'd1442,  14'd883,  14'd1123,  -14'd698,  -14'd976,  -14'd1035,  
14'd1084,  14'd2147,  -14'd860,  -14'd105,  -14'd674,  14'd1564,  14'd518,  -14'd376,  14'd983,  14'd495,  14'd1079,  -14'd762,  14'd1196,  14'd875,  -14'd373,  14'd671,  
-14'd372,  14'd1682,  14'd1789,  14'd56,  14'd1334,  14'd1626,  -14'd1551,  14'd255,  -14'd562,  14'd176,  -14'd1070,  -14'd271,  14'd1039,  14'd691,  14'd303,  14'd832,  
14'd1184,  14'd307,  14'd1395,  14'd1195,  -14'd278,  14'd967,  -14'd756,  -14'd162,  14'd1631,  -14'd172,  -14'd625,  14'd552,  -14'd347,  14'd814,  14'd109,  -14'd136,  
14'd797,  14'd709,  14'd2367,  14'd1376,  -14'd534,  14'd4,  -14'd1202,  14'd252,  -14'd395,  -14'd21,  14'd997,  -14'd626,  -14'd1531,  14'd1487,  14'd564,  -14'd469,  
14'd39,  14'd1147,  14'd2011,  -14'd1305,  -14'd696,  14'd103,  14'd135,  -14'd344,  -14'd271,  -14'd724,  -14'd827,  14'd203,  14'd372,  14'd759,  -14'd753,  -14'd541,  
14'd506,  14'd249,  -14'd1063,  14'd1125,  14'd17,  -14'd1620,  -14'd268,  -14'd383,  14'd622,  -14'd611,  14'd1648,  -14'd687,  -14'd339,  14'd226,  -14'd946,  14'd31,  
-14'd1206,  14'd331,  -14'd1077,  14'd995,  14'd780,  14'd352,  -14'd499,  14'd1202,  14'd852,  14'd561,  14'd1523,  14'd647,  14'd880,  14'd31,  14'd492,  14'd581,  
-14'd199,  -14'd801,  -14'd6,  14'd689,  14'd1324,  -14'd132,  14'd1319,  -14'd300,  14'd1239,  14'd146,  -14'd992,  -14'd834,  14'd346,  -14'd118,  14'd996,  14'd1076,  
-14'd799,  14'd645,  14'd1950,  -14'd728,  -14'd273,  14'd175,  -14'd716,  14'd885,  -14'd322,  -14'd934,  -14'd194,  14'd325,  -14'd115,  14'd963,  -14'd556,  -14'd636,  
-14'd1601,  -14'd777,  -14'd1721,  14'd1006,  -14'd199,  -14'd456,  -14'd402,  14'd878,  -14'd563,  14'd628,  14'd967,  -14'd13,  -14'd1270,  -14'd800,  14'd893,  14'd54,  
-14'd1802,  14'd163,  14'd1449,  14'd612,  -14'd59,  -14'd1244,  -14'd106,  14'd231,  -14'd971,  14'd399,  14'd1115,  -14'd1977,  -14'd588,  -14'd1538,  14'd1353,  -14'd569,  
-14'd1418,  14'd408,  -14'd470,  -14'd336,  -14'd335,  -14'd140,  -14'd481,  -14'd1385,  14'd457,  14'd439,  14'd1690,  -14'd334,  -14'd37,  -14'd1128,  -14'd742,  -14'd151,  
14'd194,  -14'd243,  14'd83,  -14'd1,  14'd706,  14'd359,  -14'd649,  -14'd77,  -14'd253,  14'd2059,  -14'd1106,  -14'd494,  -14'd462,  14'd820,  -14'd959,  -14'd170,  
-14'd1903,  14'd125,  14'd351,  -14'd292,  14'd418,  -14'd903,  -14'd1091,  14'd322,  -14'd980,  14'd432,  -14'd1805,  -14'd282,  14'd720,  14'd1409,  14'd1093,  -14'd886,  
-14'd1107,  14'd228,  14'd15,  -14'd369,  -14'd1638,  -14'd234,  14'd1117,  -14'd990,  -14'd382,  -14'd609,  14'd526,  14'd799,  -14'd1385,  -14'd1413,  -14'd314,  -14'd35,  
14'd753,  14'd802,  14'd2093,  -14'd1596,  14'd174,  14'd1201,  -14'd422,  14'd588,  -14'd401,  14'd427,  14'd960,  14'd1925,  -14'd169,  14'd305,  -14'd1069,  -14'd196,  
-14'd912,  -14'd480,  -14'd699,  -14'd1228,  -14'd435,  14'd292,  14'd214,  -14'd114,  -14'd258,  14'd763,  -14'd898,  -14'd1212,  -14'd989,  -14'd522,  -14'd334,  14'd567,  
-14'd298,  -14'd964,  14'd297,  14'd103,  -14'd345,  -14'd289,  -14'd672,  -14'd47,  -14'd892,  14'd159,  14'd302,  -14'd1188,  -14'd159,  14'd2760,  14'd1368,  14'd725,  
-14'd669,  14'd286,  14'd1475,  -14'd138,  -14'd1063,  14'd953,  -14'd673,  -14'd903,  -14'd925,  -14'd963,  -14'd1249,  -14'd130,  -14'd543,  -14'd101,  14'd478,  -14'd505,  
14'd1124,  14'd1091,  14'd364,  -14'd815,  14'd864,  -14'd1142,  -14'd75,  -14'd620,  -14'd802,  -14'd1407,  14'd2022,  -14'd632,  -14'd343,  -14'd109,  -14'd171,  14'd696,  
14'd859,  -14'd370,  -14'd549,  14'd411,  14'd1178,  14'd809,  14'd270,  -14'd478,  14'd108,  -14'd1886,  -14'd351,  14'd1231,  -14'd268,  14'd1089,  14'd504,  14'd90,  

14'd510,  14'd1638,  14'd879,  -14'd85,  -14'd495,  14'd1656,  -14'd2575,  14'd870,  14'd1295,  14'd458,  14'd435,  -14'd2011,  14'd1308,  -14'd136,  -14'd83,  14'd1266,  
-14'd493,  14'd2025,  14'd1684,  14'd413,  14'd549,  -14'd230,  -14'd11,  14'd1086,  14'd994,  -14'd1113,  14'd1310,  14'd380,  -14'd442,  14'd38,  14'd1829,  -14'd380,  
-14'd49,  14'd280,  14'd284,  -14'd387,  -14'd621,  14'd175,  -14'd195,  -14'd690,  14'd485,  -14'd1309,  14'd15,  -14'd5,  -14'd250,  14'd339,  14'd1461,  14'd1160,  
-14'd558,  -14'd404,  -14'd180,  14'd300,  -14'd1688,  14'd2270,  14'd533,  14'd949,  -14'd234,  -14'd838,  14'd1990,  14'd177,  14'd467,  14'd1189,  14'd1106,  -14'd606,  
14'd1361,  14'd287,  14'd6,  -14'd208,  -14'd1690,  14'd1068,  14'd118,  -14'd639,  -14'd125,  -14'd1480,  -14'd157,  -14'd640,  14'd336,  14'd751,  -14'd1361,  14'd86,  
-14'd1716,  14'd957,  14'd417,  -14'd2187,  14'd1887,  -14'd472,  14'd1829,  -14'd114,  -14'd99,  14'd1014,  -14'd3,  -14'd933,  14'd160,  -14'd420,  -14'd894,  -14'd283,  
-14'd1094,  -14'd801,  -14'd365,  -14'd2160,  14'd668,  14'd1670,  -14'd865,  14'd125,  -14'd491,  -14'd644,  -14'd1944,  -14'd1058,  14'd322,  14'd671,  -14'd576,  -14'd867,  
14'd449,  -14'd430,  14'd936,  -14'd344,  -14'd1734,  -14'd1612,  -14'd1416,  -14'd1311,  -14'd1494,  14'd266,  -14'd26,  -14'd54,  -14'd1246,  -14'd186,  14'd308,  -14'd804,  
-14'd289,  -14'd127,  -14'd129,  -14'd955,  -14'd1856,  14'd688,  -14'd260,  -14'd736,  -14'd62,  -14'd447,  14'd98,  -14'd1137,  -14'd1632,  14'd421,  -14'd61,  -14'd1718,  
-14'd1841,  -14'd1253,  14'd2107,  14'd121,  -14'd1199,  -14'd889,  -14'd72,  14'd698,  -14'd1261,  14'd373,  14'd155,  -14'd821,  -14'd1324,  14'd324,  14'd316,  14'd650,  
-14'd610,  -14'd909,  -14'd862,  -14'd483,  -14'd792,  -14'd711,  14'd486,  14'd578,  14'd1563,  -14'd299,  -14'd1756,  -14'd1040,  -14'd1155,  -14'd153,  14'd19,  -14'd409,  
-14'd617,  -14'd1294,  14'd91,  14'd1283,  -14'd410,  -14'd132,  14'd674,  -14'd1095,  -14'd236,  14'd84,  -14'd1850,  14'd981,  -14'd87,  -14'd170,  14'd600,  -14'd1548,  
14'd108,  -14'd127,  14'd1739,  14'd238,  14'd668,  -14'd898,  -14'd988,  -14'd288,  14'd2134,  -14'd168,  14'd143,  14'd2057,  -14'd238,  14'd2010,  -14'd1857,  14'd365,  
-14'd1553,  -14'd786,  -14'd2383,  14'd820,  -14'd112,  14'd339,  14'd435,  -14'd806,  -14'd870,  -14'd1326,  14'd1398,  14'd659,  14'd267,  14'd1030,  -14'd1468,  -14'd173,  
14'd826,  -14'd77,  14'd2451,  -14'd633,  14'd2201,  -14'd702,  -14'd1267,  -14'd797,  14'd785,  14'd873,  -14'd240,  14'd1309,  14'd1187,  14'd71,  -14'd562,  -14'd75,  
14'd1651,  14'd761,  14'd456,  -14'd1171,  -14'd2183,  14'd500,  14'd920,  -14'd1060,  14'd157,  14'd704,  -14'd625,  14'd983,  -14'd365,  14'd855,  14'd604,  14'd993,  
14'd1159,  -14'd971,  14'd1743,  14'd1464,  -14'd1550,  -14'd990,  14'd568,  14'd678,  14'd105,  -14'd1084,  14'd2061,  14'd1589,  -14'd979,  -14'd691,  14'd463,  14'd554,  
-14'd840,  14'd258,  14'd1033,  14'd1387,  14'd1626,  -14'd908,  14'd810,  -14'd1262,  14'd1738,  -14'd560,  -14'd433,  14'd602,  14'd283,  -14'd1102,  -14'd910,  -14'd552,  
-14'd420,  14'd227,  -14'd2496,  14'd89,  14'd300,  -14'd600,  14'd274,  14'd1145,  -14'd640,  14'd344,  14'd195,  14'd1733,  14'd53,  -14'd460,  14'd438,  14'd586,  
14'd693,  14'd935,  -14'd914,  -14'd1734,  -14'd3,  -14'd677,  -14'd156,  -14'd792,  14'd117,  14'd609,  -14'd1503,  -14'd496,  14'd909,  14'd1236,  14'd1730,  14'd915,  
14'd1293,  14'd574,  14'd1848,  -14'd536,  14'd1270,  -14'd120,  -14'd574,  -14'd43,  -14'd1133,  14'd152,  -14'd1414,  14'd51,  -14'd706,  14'd2253,  14'd295,  -14'd751,  
-14'd409,  14'd1716,  -14'd28,  -14'd949,  -14'd1696,  -14'd111,  14'd146,  -14'd316,  -14'd1465,  -14'd83,  14'd1203,  -14'd352,  -14'd157,  -14'd2161,  14'd1452,  -14'd86,  
-14'd1596,  14'd566,  -14'd666,  14'd734,  -14'd1187,  -14'd429,  -14'd1462,  14'd562,  14'd691,  -14'd988,  14'd989,  -14'd651,  14'd353,  14'd5,  14'd522,  -14'd1098,  
14'd866,  14'd1125,  -14'd6,  -14'd582,  -14'd136,  14'd872,  -14'd630,  -14'd1354,  14'd751,  14'd515,  14'd140,  -14'd748,  -14'd374,  14'd149,  14'd1076,  -14'd236,  
-14'd830,  14'd733,  -14'd989,  14'd1684,  14'd1130,  14'd1349,  -14'd323,  14'd633,  14'd17,  14'd437,  14'd1249,  14'd101,  14'd1474,  -14'd502,  14'd295,  14'd293,  

-14'd1241,  14'd1400,  14'd473,  14'd274,  14'd898,  -14'd183,  -14'd2236,  14'd759,  14'd46,  14'd1095,  14'd1644,  -14'd477,  -14'd230,  -14'd750,  14'd829,  -14'd33,  
-14'd1002,  -14'd954,  -14'd1332,  14'd1342,  14'd1538,  -14'd205,  -14'd496,  14'd627,  14'd428,  14'd409,  14'd1694,  -14'd108,  14'd1292,  14'd1282,  -14'd27,  14'd785,  
-14'd1736,  14'd1163,  14'd4,  14'd637,  14'd91,  14'd760,  -14'd174,  14'd695,  14'd220,  -14'd899,  -14'd12,  14'd476,  14'd731,  -14'd1557,  14'd729,  14'd1922,  
-14'd1494,  -14'd548,  -14'd1655,  14'd326,  -14'd391,  -14'd928,  -14'd1145,  14'd534,  -14'd577,  14'd234,  -14'd199,  -14'd308,  14'd1611,  -14'd805,  14'd736,  14'd805,  
14'd61,  -14'd1517,  14'd863,  14'd172,  -14'd103,  14'd939,  14'd641,  -14'd120,  -14'd1600,  -14'd788,  14'd688,  14'd275,  14'd773,  -14'd1200,  -14'd1516,  14'd724,  
-14'd189,  -14'd140,  14'd42,  14'd432,  14'd458,  14'd106,  -14'd65,  14'd1303,  -14'd1142,  14'd772,  -14'd86,  14'd928,  14'd209,  14'd158,  -14'd449,  14'd855,  
-14'd335,  -14'd1456,  -14'd611,  14'd309,  -14'd927,  -14'd261,  14'd62,  14'd1404,  -14'd1572,  14'd29,  14'd1254,  -14'd337,  14'd187,  -14'd898,  -14'd503,  -14'd407,  
-14'd1048,  14'd350,  14'd418,  -14'd254,  -14'd105,  -14'd117,  -14'd295,  14'd276,  -14'd821,  14'd547,  14'd87,  -14'd701,  -14'd691,  14'd1629,  -14'd1092,  14'd1284,  
-14'd465,  14'd1763,  14'd821,  14'd708,  -14'd236,  -14'd553,  14'd1263,  14'd513,  -14'd897,  -14'd209,  14'd80,  14'd1432,  14'd639,  14'd685,  14'd479,  -14'd170,  
14'd43,  14'd1546,  14'd506,  -14'd197,  14'd784,  -14'd490,  -14'd1247,  14'd1522,  -14'd1604,  -14'd175,  -14'd309,  -14'd341,  -14'd955,  -14'd290,  14'd757,  14'd624,  
14'd407,  -14'd109,  -14'd571,  -14'd58,  -14'd1701,  14'd242,  -14'd326,  -14'd1666,  14'd1253,  14'd260,  14'd498,  -14'd59,  -14'd1244,  -14'd1276,  -14'd1521,  -14'd474,  
14'd910,  -14'd1424,  -14'd370,  -14'd157,  -14'd369,  -14'd795,  14'd796,  14'd82,  -14'd21,  14'd196,  14'd975,  -14'd825,  14'd837,  -14'd554,  14'd91,  -14'd38,  
-14'd285,  -14'd757,  -14'd454,  14'd16,  -14'd68,  -14'd175,  14'd734,  -14'd163,  14'd937,  14'd646,  -14'd116,  -14'd646,  14'd711,  14'd982,  -14'd1226,  14'd634,  
14'd1537,  14'd760,  14'd896,  14'd311,  14'd590,  -14'd1466,  14'd157,  14'd693,  -14'd80,  -14'd1896,  -14'd888,  -14'd1053,  -14'd1422,  -14'd492,  14'd904,  -14'd1088,  
-14'd506,  14'd410,  14'd1094,  14'd498,  14'd1944,  14'd807,  -14'd69,  -14'd187,  14'd868,  -14'd351,  -14'd1154,  14'd748,  14'd1038,  14'd596,  -14'd127,  -14'd535,  
-14'd408,  -14'd112,  -14'd828,  -14'd377,  14'd744,  14'd377,  14'd262,  14'd32,  14'd1001,  14'd1080,  14'd1019,  14'd190,  14'd1028,  -14'd1078,  14'd168,  -14'd226,  
-14'd324,  -14'd644,  -14'd1112,  14'd440,  -14'd342,  14'd556,  -14'd92,  -14'd4,  14'd1002,  14'd905,  14'd146,  -14'd325,  14'd716,  14'd295,  14'd804,  -14'd722,  
14'd1057,  14'd157,  -14'd272,  14'd660,  -14'd479,  14'd797,  -14'd529,  -14'd961,  14'd422,  14'd572,  -14'd468,  14'd121,  14'd732,  14'd2452,  -14'd366,  14'd630,  
-14'd730,  -14'd447,  14'd1182,  14'd998,  14'd103,  -14'd304,  14'd282,  -14'd1157,  14'd725,  -14'd681,  14'd159,  14'd1380,  14'd348,  -14'd271,  -14'd369,  -14'd623,  
-14'd492,  -14'd1189,  14'd215,  14'd576,  14'd1691,  -14'd628,  -14'd445,  14'd221,  14'd534,  14'd1185,  -14'd117,  14'd1015,  14'd1084,  14'd316,  14'd178,  -14'd1060,  
14'd57,  -14'd171,  14'd190,  -14'd920,  -14'd1889,  -14'd513,  14'd1140,  14'd56,  14'd287,  -14'd544,  14'd1599,  -14'd1278,  -14'd709,  14'd854,  -14'd439,  -14'd128,  
14'd49,  14'd400,  -14'd564,  14'd1189,  -14'd665,  14'd1076,  14'd1838,  14'd1760,  14'd541,  14'd443,  14'd1339,  -14'd472,  14'd169,  14'd1005,  14'd1965,  14'd78,  
-14'd406,  -14'd1122,  14'd883,  14'd716,  -14'd916,  -14'd1255,  -14'd774,  -14'd778,  -14'd1112,  -14'd909,  -14'd1411,  -14'd727,  -14'd984,  14'd2029,  14'd1044,  14'd681,  
-14'd1415,  14'd401,  -14'd417,  -14'd210,  14'd70,  -14'd285,  14'd604,  -14'd254,  -14'd72,  -14'd462,  -14'd250,  -14'd417,  14'd714,  -14'd591,  14'd537,  14'd662,  
14'd77,  14'd2204,  -14'd172,  14'd355,  14'd1536,  14'd1135,  -14'd1213,  -14'd675,  14'd341,  14'd1322,  14'd255,  -14'd210,  -14'd457,  14'd786,  -14'd1197,  14'd351,  

-14'd1522,  -14'd57,  -14'd203,  -14'd230,  -14'd857,  14'd636,  14'd1402,  14'd699,  -14'd1141,  14'd278,  14'd505,  14'd204,  14'd497,  14'd1077,  14'd242,  -14'd851,  
14'd1417,  -14'd176,  14'd88,  -14'd130,  14'd808,  14'd688,  14'd1284,  14'd707,  -14'd881,  14'd600,  14'd2093,  14'd1315,  -14'd267,  14'd465,  14'd405,  14'd454,  
14'd642,  14'd225,  -14'd158,  14'd1164,  14'd1509,  14'd528,  14'd886,  14'd152,  14'd529,  -14'd242,  14'd1285,  14'd535,  -14'd153,  14'd1046,  14'd966,  -14'd684,  
-14'd81,  14'd2261,  14'd1442,  -14'd116,  -14'd296,  14'd190,  -14'd1025,  14'd375,  14'd317,  -14'd488,  -14'd539,  14'd940,  14'd555,  -14'd949,  -14'd1145,  14'd1413,  
-14'd213,  14'd368,  14'd696,  -14'd290,  -14'd131,  14'd4,  -14'd1723,  14'd394,  14'd948,  14'd624,  14'd67,  14'd61,  -14'd124,  14'd800,  -14'd778,  -14'd455,  
14'd546,  -14'd377,  -14'd1301,  -14'd47,  -14'd79,  -14'd1633,  14'd31,  14'd21,  -14'd1057,  -14'd234,  14'd1208,  -14'd893,  14'd18,  14'd293,  -14'd960,  -14'd193,  
-14'd790,  -14'd194,  14'd2023,  14'd866,  -14'd829,  14'd1403,  14'd2203,  -14'd843,  14'd83,  14'd323,  -14'd630,  -14'd101,  -14'd1419,  14'd283,  14'd406,  -14'd840,  
-14'd1445,  14'd1881,  14'd46,  14'd140,  14'd1268,  -14'd105,  14'd1052,  -14'd578,  14'd1056,  14'd571,  14'd1137,  -14'd2013,  -14'd349,  -14'd75,  -14'd570,  -14'd891,  
-14'd2305,  -14'd71,  -14'd959,  -14'd978,  14'd1457,  -14'd613,  -14'd2049,  -14'd643,  -14'd282,  14'd1563,  -14'd556,  -14'd673,  -14'd1487,  -14'd791,  14'd255,  -14'd121,  
-14'd4140,  -14'd1934,  14'd1347,  -14'd1296,  -14'd1562,  14'd8,  -14'd1246,  -14'd354,  -14'd847,  -14'd433,  -14'd73,  -14'd1515,  -14'd1973,  -14'd115,  14'd1825,  14'd237,  
-14'd81,  -14'd1127,  -14'd651,  -14'd570,  -14'd1363,  -14'd838,  14'd2579,  -14'd896,  14'd662,  -14'd917,  -14'd83,  14'd665,  -14'd810,  -14'd620,  14'd31,  14'd457,  
14'd1394,  -14'd1212,  14'd184,  14'd120,  -14'd1403,  -14'd808,  -14'd1389,  14'd376,  14'd137,  14'd119,  -14'd977,  -14'd921,  -14'd267,  -14'd475,  -14'd1465,  -14'd398,  
-14'd1699,  -14'd114,  -14'd49,  -14'd227,  14'd532,  -14'd1664,  -14'd1193,  14'd456,  14'd1052,  14'd953,  -14'd1706,  -14'd280,  -14'd1632,  14'd340,  -14'd140,  -14'd556,  
-14'd484,  14'd941,  14'd568,  -14'd140,  -14'd880,  14'd406,  14'd190,  -14'd2014,  14'd1140,  -14'd899,  -14'd1475,  14'd319,  -14'd858,  14'd1186,  -14'd491,  -14'd1827,  
-14'd635,  -14'd286,  14'd2051,  14'd129,  -14'd592,  -14'd234,  -14'd159,  -14'd137,  14'd1097,  14'd130,  -14'd1542,  14'd2397,  -14'd1502,  14'd1246,  14'd988,  -14'd2234,  
14'd1716,  14'd711,  14'd786,  -14'd354,  -14'd1625,  14'd516,  14'd46,  14'd716,  14'd88,  14'd1311,  -14'd1626,  14'd103,  14'd1485,  14'd705,  14'd398,  14'd128,  
-14'd333,  -14'd18,  14'd457,  -14'd597,  -14'd1200,  14'd898,  14'd571,  14'd1001,  14'd715,  -14'd240,  14'd921,  14'd811,  -14'd770,  14'd2322,  14'd1162,  14'd1813,  
14'd465,  -14'd1587,  14'd551,  14'd782,  -14'd728,  14'd601,  -14'd356,  14'd536,  -14'd473,  14'd253,  14'd344,  14'd657,  14'd111,  14'd522,  -14'd504,  14'd1373,  
14'd99,  14'd803,  14'd1153,  14'd1229,  -14'd336,  -14'd103,  14'd313,  -14'd818,  14'd347,  -14'd545,  -14'd186,  14'd101,  14'd1070,  14'd775,  14'd529,  -14'd529,  
14'd2679,  -14'd11,  14'd974,  14'd1618,  14'd618,  -14'd603,  14'd330,  -14'd94,  -14'd1214,  14'd1004,  14'd652,  14'd1425,  14'd1532,  -14'd1494,  14'd161,  -14'd1209,  
-14'd271,  -14'd246,  -14'd608,  14'd383,  -14'd597,  -14'd863,  -14'd46,  -14'd455,  -14'd1023,  -14'd213,  -14'd822,  -14'd112,  -14'd437,  14'd69,  -14'd127,  14'd372,  
-14'd869,  14'd672,  -14'd351,  14'd1193,  14'd20,  14'd124,  14'd848,  -14'd1238,  -14'd347,  14'd136,  14'd333,  -14'd371,  -14'd172,  14'd1651,  14'd834,  14'd152,  
-14'd75,  14'd957,  14'd943,  14'd416,  -14'd298,  14'd443,  14'd831,  14'd473,  14'd485,  14'd437,  -14'd23,  -14'd617,  -14'd311,  -14'd963,  -14'd717,  14'd218,  
-14'd294,  14'd1614,  -14'd577,  -14'd331,  14'd66,  -14'd640,  -14'd1004,  14'd239,  14'd129,  -14'd1265,  -14'd3,  -14'd1669,  14'd835,  -14'd944,  -14'd311,  14'd1439,  
-14'd475,  14'd949,  -14'd1737,  -14'd306,  14'd710,  -14'd636,  -14'd246,  14'd680,  -14'd899,  14'd40,  -14'd781,  -14'd324,  -14'd274,  -14'd262,  -14'd420,  14'd124,  

-14'd289,  14'd1512,  -14'd513,  -14'd314,  14'd238,  -14'd106,  -14'd678,  -14'd202,  14'd549,  14'd226,  -14'd650,  -14'd333,  14'd1426,  -14'd1207,  14'd370,  14'd562,  
-14'd550,  -14'd366,  -14'd1526,  14'd188,  14'd452,  14'd932,  -14'd991,  14'd277,  -14'd264,  -14'd707,  -14'd1253,  14'd368,  14'd1037,  -14'd339,  14'd1143,  14'd892,  
-14'd545,  -14'd796,  14'd630,  14'd557,  -14'd553,  -14'd557,  14'd1320,  14'd112,  -14'd1462,  -14'd50,  14'd836,  -14'd325,  14'd711,  -14'd2042,  14'd102,  14'd389,  
-14'd769,  -14'd589,  -14'd581,  -14'd433,  -14'd606,  14'd730,  14'd1545,  -14'd1117,  14'd757,  -14'd64,  14'd1169,  14'd694,  -14'd1429,  14'd943,  -14'd952,  14'd398,  
-14'd379,  14'd1062,  -14'd960,  14'd48,  -14'd639,  -14'd485,  14'd1036,  14'd40,  -14'd665,  -14'd825,  14'd36,  -14'd82,  -14'd1181,  14'd130,  -14'd1671,  14'd109,  
14'd429,  14'd202,  14'd49,  14'd1387,  -14'd99,  -14'd359,  -14'd1115,  14'd1225,  -14'd872,  -14'd2293,  14'd838,  14'd198,  -14'd749,  14'd741,  -14'd220,  14'd672,  
-14'd1136,  14'd507,  14'd30,  -14'd329,  14'd243,  14'd1176,  -14'd277,  -14'd133,  -14'd997,  14'd387,  14'd1060,  -14'd119,  14'd1052,  -14'd1741,  14'd1062,  14'd1290,  
-14'd370,  14'd4,  -14'd1347,  -14'd1089,  14'd1522,  -14'd973,  14'd296,  -14'd219,  14'd425,  -14'd530,  14'd1202,  14'd112,  -14'd687,  -14'd848,  -14'd114,  14'd1601,  
14'd264,  -14'd439,  -14'd666,  -14'd976,  -14'd606,  14'd689,  14'd992,  14'd369,  14'd872,  14'd861,  14'd262,  -14'd647,  -14'd61,  14'd592,  -14'd289,  -14'd525,  
14'd1047,  14'd1373,  14'd1258,  14'd899,  14'd35,  -14'd600,  -14'd1044,  14'd610,  -14'd104,  14'd1304,  14'd156,  -14'd1496,  14'd1135,  14'd536,  -14'd366,  -14'd537,  
14'd971,  14'd36,  14'd664,  -14'd728,  -14'd1375,  -14'd782,  -14'd973,  14'd543,  14'd626,  14'd234,  14'd756,  -14'd1326,  14'd1284,  14'd417,  14'd132,  -14'd424,  
-14'd349,  14'd673,  -14'd425,  14'd42,  14'd863,  -14'd128,  -14'd1723,  -14'd46,  -14'd997,  14'd291,  14'd150,  14'd831,  14'd629,  -14'd768,  -14'd687,  14'd281,  
-14'd1266,  -14'd875,  14'd1375,  -14'd776,  -14'd166,  14'd1163,  -14'd778,  -14'd107,  -14'd1507,  -14'd308,  -14'd538,  14'd78,  14'd919,  -14'd51,  14'd932,  -14'd844,  
-14'd655,  -14'd979,  -14'd1390,  14'd627,  14'd784,  14'd293,  14'd9,  -14'd1613,  14'd167,  14'd973,  -14'd429,  -14'd566,  14'd425,  -14'd1681,  14'd62,  14'd543,  
-14'd1918,  -14'd921,  14'd939,  14'd804,  -14'd118,  -14'd52,  -14'd1204,  -14'd9,  14'd836,  14'd2325,  -14'd15,  14'd625,  -14'd979,  14'd1358,  -14'd965,  -14'd961,  
-14'd1793,  14'd407,  -14'd95,  14'd39,  -14'd197,  -14'd45,  -14'd868,  -14'd492,  14'd2418,  -14'd64,  14'd992,  -14'd2044,  -14'd993,  -14'd1595,  -14'd831,  -14'd1664,  
-14'd1023,  -14'd543,  -14'd1169,  -14'd640,  -14'd1008,  14'd370,  -14'd836,  -14'd675,  -14'd517,  14'd1649,  14'd1336,  -14'd1281,  14'd468,  -14'd1318,  -14'd1250,  -14'd893,  
-14'd88,  -14'd296,  14'd668,  -14'd322,  14'd374,  -14'd644,  -14'd494,  -14'd91,  -14'd555,  -14'd265,  14'd157,  -14'd327,  -14'd541,  -14'd1106,  -14'd373,  14'd657,  
-14'd467,  -14'd13,  -14'd853,  14'd944,  14'd1585,  14'd1001,  -14'd1362,  14'd110,  -14'd747,  -14'd1053,  -14'd692,  14'd1044,  14'd1578,  -14'd1111,  -14'd263,  14'd365,  
-14'd1424,  -14'd271,  14'd289,  14'd1196,  -14'd152,  14'd689,  14'd477,  -14'd452,  14'd669,  14'd856,  -14'd205,  14'd556,  14'd162,  14'd338,  -14'd1008,  -14'd1213,  
-14'd297,  -14'd362,  -14'd1241,  14'd1020,  14'd429,  14'd681,  14'd2258,  -14'd880,  14'd1215,  14'd378,  14'd1770,  -14'd861,  -14'd458,  -14'd614,  -14'd131,  -14'd1017,  
14'd1247,  14'd168,  -14'd256,  -14'd193,  -14'd940,  -14'd1319,  14'd69,  -14'd1143,  14'd2224,  14'd1590,  -14'd177,  14'd885,  14'd649,  -14'd2281,  -14'd441,  14'd78,  
14'd570,  14'd1110,  -14'd683,  14'd901,  14'd12,  14'd76,  -14'd509,  -14'd112,  14'd1533,  14'd2005,  14'd868,  14'd1230,  -14'd709,  14'd361,  -14'd805,  14'd1060,  
14'd1610,  14'd1102,  -14'd1047,  -14'd851,  14'd1006,  14'd1205,  -14'd472,  14'd763,  14'd700,  -14'd838,  -14'd106,  -14'd901,  14'd1523,  14'd1298,  -14'd242,  -14'd600,  
14'd402,  14'd325,  14'd1497,  14'd407,  -14'd194,  14'd743,  -14'd619,  -14'd959,  14'd1426,  14'd249,  -14'd380,  -14'd984,  -14'd218,  14'd1063,  -14'd1141,  14'd723,  

14'd1745,  -14'd1753,  -14'd971,  14'd113,  -14'd1530,  14'd885,  14'd384,  -14'd546,  -14'd1030,  14'd587,  14'd1242,  14'd215,  -14'd759,  14'd845,  -14'd1584,  -14'd740,  
-14'd407,  -14'd687,  -14'd129,  -14'd1302,  -14'd1113,  14'd356,  14'd250,  -14'd2104,  14'd120,  -14'd241,  -14'd279,  14'd1525,  -14'd321,  14'd503,  14'd330,  14'd143,  
14'd699,  14'd3,  -14'd172,  -14'd569,  14'd661,  -14'd533,  -14'd1314,  14'd1166,  14'd1432,  -14'd301,  -14'd374,  14'd735,  14'd558,  -14'd373,  -14'd303,  14'd1238,  
-14'd84,  14'd339,  -14'd417,  14'd520,  -14'd526,  -14'd164,  14'd317,  14'd441,  14'd739,  -14'd737,  -14'd1541,  -14'd725,  -14'd1197,  14'd496,  14'd658,  14'd758,  
-14'd1170,  14'd325,  -14'd2,  14'd166,  14'd171,  -14'd268,  14'd1078,  14'd50,  14'd572,  -14'd111,  -14'd1242,  14'd358,  14'd2,  14'd719,  -14'd1303,  -14'd921,  
14'd204,  -14'd305,  14'd425,  14'd699,  14'd383,  14'd780,  14'd1757,  -14'd936,  14'd1497,  -14'd590,  14'd403,  14'd1442,  -14'd84,  14'd770,  -14'd937,  -14'd1112,  
14'd262,  14'd566,  14'd321,  14'd671,  -14'd13,  -14'd208,  14'd938,  -14'd1154,  14'd1972,  14'd845,  -14'd1919,  14'd240,  -14'd312,  14'd1044,  14'd1283,  14'd1133,  
14'd1364,  14'd1133,  14'd152,  -14'd48,  14'd1025,  -14'd262,  14'd1262,  14'd180,  -14'd1072,  -14'd582,  -14'd397,  14'd641,  -14'd711,  -14'd249,  14'd364,  -14'd12,  
-14'd968,  -14'd781,  14'd48,  14'd143,  14'd1037,  -14'd651,  14'd27,  -14'd1509,  14'd797,  -14'd475,  -14'd1550,  14'd872,  -14'd20,  14'd764,  -14'd876,  14'd839,  
14'd1635,  -14'd473,  -14'd1354,  14'd1288,  -14'd640,  -14'd1318,  14'd1087,  -14'd600,  14'd17,  -14'd1450,  14'd741,  14'd510,  14'd467,  -14'd144,  14'd575,  14'd847,  
14'd738,  14'd446,  14'd2008,  14'd173,  14'd520,  14'd312,  14'd1035,  14'd826,  -14'd793,  14'd415,  -14'd1915,  14'd1496,  14'd313,  14'd536,  14'd141,  14'd1237,  
14'd620,  14'd203,  14'd176,  14'd193,  14'd1486,  -14'd110,  14'd220,  14'd747,  14'd405,  14'd307,  -14'd840,  14'd413,  14'd350,  14'd247,  -14'd997,  -14'd252,  
14'd704,  -14'd129,  -14'd290,  14'd475,  -14'd1748,  14'd978,  14'd986,  14'd174,  -14'd1106,  -14'd1448,  -14'd642,  14'd431,  -14'd1609,  -14'd731,  -14'd607,  14'd644,  
14'd727,  -14'd121,  -14'd1156,  -14'd105,  -14'd1273,  14'd726,  14'd87,  14'd112,  14'd226,  -14'd491,  14'd7,  14'd372,  14'd763,  14'd988,  -14'd368,  -14'd691,  
-14'd10,  -14'd16,  -14'd1069,  -14'd9,  14'd1212,  14'd934,  -14'd50,  -14'd617,  -14'd1164,  -14'd377,  14'd63,  -14'd426,  14'd1763,  -14'd53,  -14'd835,  14'd810,  
14'd947,  14'd458,  14'd1390,  14'd124,  14'd777,  -14'd62,  14'd288,  14'd683,  -14'd1268,  14'd781,  -14'd1913,  14'd1622,  14'd988,  14'd650,  14'd680,  14'd14,  
14'd698,  14'd1203,  -14'd43,  -14'd1225,  -14'd324,  14'd65,  14'd247,  -14'd0,  -14'd1090,  14'd171,  -14'd963,  -14'd1528,  14'd1362,  14'd291,  -14'd214,  14'd935,  
14'd1434,  -14'd42,  -14'd695,  -14'd466,  -14'd915,  -14'd1032,  14'd108,  14'd1154,  -14'd689,  -14'd453,  14'd32,  -14'd908,  -14'd1444,  14'd720,  -14'd530,  14'd465,  
14'd70,  14'd103,  -14'd406,  -14'd920,  14'd1233,  -14'd1832,  14'd1217,  -14'd156,  -14'd772,  -14'd62,  14'd111,  -14'd588,  -14'd1255,  -14'd1383,  14'd301,  14'd691,  
-14'd1348,  -14'd920,  -14'd412,  14'd1259,  -14'd489,  -14'd898,  -14'd492,  -14'd800,  14'd155,  -14'd612,  14'd626,  14'd159,  -14'd1355,  -14'd320,  -14'd774,  14'd263,  
14'd1019,  14'd164,  14'd195,  14'd1321,  -14'd614,  14'd1037,  -14'd1037,  14'd343,  -14'd2646,  14'd1472,  -14'd1065,  -14'd109,  -14'd564,  14'd2023,  14'd222,  -14'd152,  
14'd538,  -14'd1076,  14'd867,  -14'd359,  -14'd1306,  -14'd1046,  -14'd802,  14'd1222,  14'd109,  14'd84,  -14'd1004,  -14'd530,  14'd614,  14'd1352,  -14'd785,  -14'd262,  
-14'd661,  14'd392,  14'd16,  14'd507,  -14'd16,  14'd180,  -14'd1751,  14'd980,  -14'd487,  -14'd933,  -14'd1096,  -14'd583,  14'd864,  14'd428,  14'd1457,  -14'd811,  
14'd104,  -14'd654,  14'd648,  14'd603,  14'd1107,  -14'd872,  -14'd537,  -14'd465,  -14'd1634,  -14'd974,  14'd127,  -14'd996,  -14'd803,  -14'd1091,  14'd994,  -14'd662,  
-14'd418,  -14'd401,  -14'd492,  14'd216,  14'd259,  14'd1089,  14'd279,  14'd359,  -14'd1071,  -14'd1922,  14'd280,  14'd862,  -14'd170,  -14'd365,  14'd1085,  -14'd431,  

-14'd1464,  -14'd846,  14'd136,  -14'd622,  -14'd1447,  -14'd436,  14'd1116,  14'd544,  14'd826,  -14'd372,  -14'd1300,  -14'd543,  -14'd2122,  -14'd95,  -14'd495,  -14'd1903,  
-14'd1022,  14'd239,  -14'd1634,  14'd1047,  14'd74,  -14'd68,  14'd167,  14'd453,  14'd1055,  -14'd880,  -14'd467,  -14'd721,  -14'd772,  -14'd65,  14'd938,  -14'd555,  
14'd345,  -14'd981,  14'd656,  -14'd830,  -14'd814,  -14'd399,  -14'd2023,  -14'd450,  14'd940,  14'd151,  -14'd424,  -14'd467,  14'd226,  -14'd876,  -14'd668,  14'd182,  
-14'd1267,  -14'd173,  -14'd478,  14'd311,  14'd756,  -14'd1480,  -14'd483,  14'd1154,  -14'd1407,  14'd981,  -14'd1064,  14'd27,  14'd1533,  -14'd2194,  14'd192,  14'd1301,  
-14'd1123,  -14'd2184,  14'd625,  -14'd285,  14'd1096,  14'd210,  -14'd45,  -14'd248,  14'd276,  -14'd1403,  14'd41,  -14'd516,  -14'd42,  14'd1433,  14'd974,  14'd269,  
-14'd426,  -14'd761,  -14'd1565,  -14'd336,  14'd345,  -14'd954,  14'd327,  -14'd64,  -14'd166,  -14'd289,  -14'd279,  -14'd380,  -14'd554,  14'd21,  -14'd1838,  -14'd956,  
-14'd473,  14'd202,  -14'd287,  -14'd683,  -14'd89,  -14'd861,  -14'd2197,  -14'd614,  -14'd1278,  14'd1822,  14'd22,  14'd661,  -14'd1336,  14'd670,  -14'd1548,  14'd1464,  
-14'd248,  -14'd449,  -14'd772,  -14'd1275,  14'd671,  14'd1038,  -14'd372,  14'd963,  14'd1103,  14'd596,  -14'd817,  14'd1586,  14'd224,  14'd53,  14'd1410,  -14'd967,  
-14'd874,  -14'd1903,  -14'd1106,  14'd390,  -14'd747,  14'd776,  -14'd645,  -14'd230,  -14'd474,  -14'd488,  14'd332,  14'd48,  -14'd301,  -14'd1031,  14'd135,  14'd962,  
-14'd191,  -14'd199,  14'd1088,  14'd921,  14'd746,  14'd635,  14'd726,  14'd1061,  -14'd1409,  -14'd367,  14'd1450,  14'd1487,  14'd1837,  -14'd1150,  -14'd41,  14'd930,  
14'd527,  14'd205,  -14'd1110,  14'd1132,  14'd210,  14'd849,  -14'd105,  14'd223,  14'd1050,  -14'd1294,  -14'd2468,  14'd68,  14'd925,  -14'd937,  -14'd165,  -14'd1096,  
-14'd1312,  14'd762,  14'd1022,  -14'd1001,  -14'd380,  14'd669,  14'd497,  -14'd1357,  14'd924,  14'd361,  14'd301,  14'd545,  -14'd295,  -14'd730,  14'd869,  -14'd1325,  
14'd554,  14'd409,  14'd721,  -14'd783,  14'd93,  -14'd496,  -14'd636,  -14'd1908,  -14'd992,  14'd1797,  14'd1568,  14'd709,  -14'd81,  14'd14,  -14'd101,  14'd579,  
14'd800,  14'd83,  14'd1019,  14'd77,  -14'd251,  -14'd1125,  14'd365,  14'd1480,  -14'd79,  14'd611,  14'd873,  -14'd742,  -14'd42,  14'd1517,  -14'd1184,  14'd832,  
-14'd385,  -14'd704,  -14'd2072,  -14'd1007,  14'd838,  -14'd477,  -14'd463,  -14'd8,  -14'd1671,  -14'd359,  14'd176,  -14'd1340,  14'd488,  14'd365,  14'd981,  14'd1312,  
14'd1061,  -14'd263,  14'd597,  14'd751,  14'd767,  14'd1611,  -14'd1251,  -14'd457,  14'd1756,  -14'd224,  -14'd654,  -14'd797,  -14'd1188,  -14'd161,  14'd931,  -14'd751,  
-14'd937,  14'd848,  14'd576,  -14'd15,  14'd384,  14'd686,  -14'd1090,  -14'd925,  14'd1865,  14'd639,  14'd440,  -14'd1441,  -14'd656,  -14'd711,  -14'd49,  14'd290,  
14'd1008,  -14'd467,  -14'd243,  14'd475,  14'd1660,  -14'd75,  14'd473,  14'd835,  -14'd247,  -14'd601,  14'd123,  14'd528,  -14'd277,  -14'd39,  14'd75,  14'd822,  
-14'd863,  -14'd313,  -14'd512,  -14'd708,  14'd631,  -14'd1114,  14'd1424,  -14'd1368,  14'd681,  14'd766,  -14'd55,  14'd295,  -14'd191,  14'd130,  14'd352,  -14'd709,  
-14'd884,  -14'd1730,  -14'd241,  -14'd916,  -14'd1840,  -14'd270,  -14'd881,  -14'd149,  -14'd1619,  -14'd1974,  -14'd1243,  -14'd210,  -14'd1536,  14'd205,  -14'd999,  -14'd994,  
-14'd341,  -14'd459,  14'd641,  14'd627,  14'd1996,  14'd672,  -14'd258,  14'd670,  14'd347,  -14'd692,  14'd1046,  -14'd367,  14'd1272,  -14'd314,  -14'd220,  -14'd896,  
14'd59,  14'd30,  14'd700,  14'd259,  14'd1142,  -14'd265,  -14'd1123,  14'd167,  -14'd1385,  -14'd931,  14'd62,  -14'd370,  14'd284,  -14'd1986,  14'd637,  -14'd577,  
14'd795,  -14'd767,  14'd872,  14'd641,  -14'd1769,  14'd1279,  14'd752,  -14'd1053,  -14'd577,  -14'd1854,  14'd517,  -14'd37,  -14'd311,  -14'd395,  -14'd745,  -14'd521,  
-14'd106,  -14'd924,  14'd102,  14'd1390,  -14'd1314,  14'd1387,  14'd1133,  -14'd1787,  14'd1698,  -14'd2475,  -14'd627,  14'd1203,  -14'd1762,  14'd411,  -14'd1111,  -14'd721,  
14'd334,  -14'd376,  14'd3221,  14'd264,  -14'd854,  14'd78,  -14'd78,  -14'd939,  14'd2835,  14'd1479,  -14'd86,  -14'd1216,  -14'd1332,  14'd1213,  -14'd2670,  -14'd1329,  

14'd148,  14'd486,  -14'd1340,  14'd576,  -14'd1073,  14'd178,  14'd1297,  14'd552,  14'd575,  14'd344,  -14'd712,  -14'd628,  14'd108,  14'd694,  14'd117,  14'd649,  
14'd753,  -14'd832,  -14'd719,  -14'd567,  -14'd129,  14'd22,  14'd1095,  -14'd990,  14'd1778,  14'd496,  -14'd1534,  -14'd430,  14'd329,  14'd1053,  14'd1626,  -14'd69,  
-14'd950,  -14'd132,  14'd15,  -14'd1144,  14'd73,  -14'd874,  14'd842,  -14'd578,  -14'd1124,  14'd710,  14'd154,  14'd598,  -14'd461,  -14'd188,  -14'd963,  14'd686,  
-14'd509,  14'd755,  14'd560,  -14'd109,  -14'd372,  -14'd1539,  14'd856,  -14'd557,  14'd833,  -14'd1324,  14'd253,  14'd575,  14'd479,  -14'd27,  -14'd855,  14'd1493,  
14'd455,  14'd2077,  -14'd913,  14'd1160,  14'd1155,  14'd72,  14'd117,  14'd833,  -14'd752,  14'd207,  14'd268,  14'd177,  14'd206,  -14'd682,  14'd897,  14'd1176,  
-14'd913,  14'd1278,  14'd288,  14'd196,  14'd19,  -14'd933,  14'd888,  14'd391,  -14'd437,  14'd1420,  -14'd416,  -14'd1631,  14'd663,  14'd675,  14'd904,  -14'd370,  
-14'd435,  -14'd1651,  -14'd29,  14'd366,  14'd882,  14'd319,  -14'd1373,  14'd64,  -14'd2234,  14'd1309,  -14'd553,  -14'd617,  14'd454,  14'd2416,  14'd1159,  -14'd755,  
14'd389,  -14'd658,  -14'd55,  14'd1373,  14'd644,  -14'd316,  14'd1062,  14'd1785,  -14'd841,  -14'd1508,  -14'd665,  14'd1002,  -14'd255,  -14'd636,  14'd1257,  14'd549,  
14'd91,  -14'd960,  14'd626,  14'd47,  -14'd417,  14'd49,  14'd1087,  14'd1079,  14'd1383,  -14'd1918,  14'd1437,  14'd470,  -14'd231,  -14'd1520,  14'd0,  -14'd1451,  
14'd2215,  -14'd1020,  -14'd1901,  -14'd1119,  14'd368,  14'd1087,  14'd379,  14'd989,  -14'd732,  -14'd1209,  14'd428,  -14'd1465,  14'd903,  14'd290,  -14'd2339,  14'd383,  
-14'd1230,  14'd579,  -14'd2042,  14'd861,  14'd1673,  -14'd290,  -14'd848,  -14'd229,  -14'd69,  -14'd1257,  -14'd924,  -14'd916,  14'd1347,  -14'd1565,  -14'd1010,  -14'd1176,  
-14'd701,  14'd1267,  -14'd432,  14'd957,  14'd160,  14'd421,  -14'd1793,  14'd474,  -14'd345,  14'd454,  -14'd99,  -14'd209,  -14'd762,  14'd1588,  14'd766,  14'd859,  
14'd1805,  14'd1481,  -14'd571,  14'd620,  14'd481,  14'd686,  -14'd472,  -14'd42,  14'd129,  14'd1192,  14'd510,  -14'd875,  14'd1059,  -14'd1408,  14'd418,  -14'd524,  
-14'd2229,  -14'd1694,  -14'd1150,  -14'd1501,  14'd90,  -14'd1532,  -14'd132,  -14'd77,  -14'd25,  -14'd301,  -14'd1564,  -14'd1933,  14'd1029,  -14'd970,  -14'd774,  14'd103,  
-14'd1564,  -14'd666,  -14'd1287,  -14'd460,  -14'd155,  14'd53,  -14'd1132,  14'd446,  -14'd1248,  14'd828,  14'd900,  -14'd160,  -14'd1211,  14'd172,  -14'd559,  14'd1621,  
-14'd860,  -14'd996,  -14'd1133,  14'd657,  14'd384,  -14'd334,  -14'd1363,  -14'd1351,  14'd287,  14'd759,  -14'd2011,  14'd675,  -14'd278,  14'd478,  -14'd50,  14'd656,  
14'd781,  14'd1349,  14'd1727,  14'd378,  14'd1667,  -14'd424,  14'd991,  -14'd393,  -14'd795,  14'd1058,  -14'd997,  -14'd70,  -14'd95,  14'd693,  -14'd850,  14'd204,  
14'd621,  14'd1023,  14'd706,  -14'd669,  14'd576,  14'd258,  14'd107,  -14'd1237,  -14'd1539,  -14'd95,  -14'd1725,  14'd885,  14'd478,  -14'd1650,  14'd184,  14'd435,  
14'd111,  -14'd1203,  -14'd724,  14'd82,  14'd1452,  14'd1040,  14'd200,  -14'd682,  14'd651,  -14'd410,  -14'd1050,  14'd1150,  14'd196,  14'd1113,  -14'd731,  -14'd540,  
-14'd630,  -14'd10,  14'd2743,  -14'd791,  -14'd1348,  -14'd21,  -14'd424,  -14'd302,  14'd165,  -14'd1673,  -14'd341,  14'd620,  14'd38,  14'd1061,  -14'd2346,  -14'd1402,  
-14'd325,  -14'd243,  14'd181,  -14'd48,  14'd1366,  -14'd40,  -14'd2255,  14'd479,  14'd2486,  -14'd1097,  -14'd199,  -14'd184,  -14'd36,  -14'd2181,  14'd39,  -14'd189,  
14'd100,  -14'd408,  -14'd460,  14'd651,  14'd1178,  14'd737,  -14'd743,  -14'd13,  14'd639,  14'd19,  14'd777,  14'd589,  14'd238,  -14'd2024,  -14'd1218,  14'd1056,  
14'd1347,  14'd759,  -14'd26,  -14'd726,  14'd564,  14'd163,  -14'd681,  -14'd19,  14'd51,  14'd1588,  14'd849,  14'd1931,  14'd1229,  -14'd993,  -14'd1185,  -14'd1276,  
14'd314,  14'd387,  14'd1147,  -14'd234,  -14'd898,  14'd1547,  14'd1105,  14'd385,  14'd1544,  14'd809,  14'd1161,  14'd1596,  14'd929,  14'd1457,  -14'd550,  -14'd556,  
14'd189,  14'd306,  14'd516,  -14'd1215,  14'd232,  14'd853,  14'd1031,  14'd1008,  14'd2368,  -14'd2392,  14'd321,  14'd645,  14'd1084,  14'd1929,  -14'd1614,  -14'd37,  

-14'd744,  14'd175,  -14'd1292,  -14'd1586,  -14'd1317,  -14'd872,  14'd667,  -14'd420,  -14'd413,  -14'd740,  14'd382,  -14'd41,  -14'd625,  -14'd1170,  -14'd721,  -14'd70,  
-14'd345,  14'd1276,  14'd338,  -14'd286,  -14'd825,  -14'd633,  -14'd311,  -14'd282,  14'd587,  14'd262,  -14'd666,  -14'd1072,  14'd7,  14'd678,  14'd700,  14'd192,  
-14'd577,  14'd1154,  14'd878,  14'd494,  -14'd1137,  14'd595,  14'd702,  14'd1059,  -14'd1232,  14'd803,  -14'd1010,  -14'd1121,  14'd482,  -14'd1892,  -14'd476,  14'd879,  
-14'd816,  -14'd1255,  14'd958,  14'd229,  14'd506,  14'd587,  -14'd683,  14'd173,  -14'd1020,  -14'd299,  -14'd672,  14'd11,  -14'd478,  14'd751,  14'd352,  -14'd111,  
-14'd1085,  -14'd26,  -14'd1076,  -14'd179,  -14'd507,  -14'd587,  14'd22,  -14'd102,  14'd264,  14'd546,  14'd738,  -14'd1382,  -14'd1309,  14'd906,  -14'd577,  -14'd623,  
-14'd1058,  14'd1027,  14'd654,  14'd429,  -14'd1120,  -14'd890,  14'd226,  -14'd663,  -14'd198,  -14'd2220,  14'd1641,  14'd969,  -14'd1031,  14'd489,  14'd767,  -14'd1224,  
14'd1991,  14'd955,  14'd937,  14'd946,  -14'd372,  -14'd855,  14'd875,  14'd203,  14'd534,  -14'd805,  -14'd1531,  -14'd104,  -14'd482,  14'd600,  14'd428,  -14'd952,  
14'd474,  -14'd713,  -14'd315,  -14'd432,  14'd202,  -14'd851,  -14'd756,  14'd537,  -14'd511,  -14'd763,  -14'd980,  14'd46,  14'd50,  -14'd1463,  14'd446,  -14'd288,  
14'd603,  14'd201,  14'd20,  14'd504,  -14'd409,  -14'd879,  14'd174,  -14'd539,  -14'd1172,  -14'd881,  -14'd183,  -14'd410,  -14'd590,  14'd613,  14'd733,  14'd1364,  
-14'd643,  14'd1645,  14'd1722,  -14'd94,  -14'd688,  14'd165,  14'd353,  14'd1823,  -14'd349,  14'd121,  -14'd892,  14'd81,  14'd356,  14'd426,  -14'd1172,  14'd724,  
14'd831,  14'd144,  14'd795,  -14'd949,  -14'd1576,  -14'd1566,  14'd2209,  -14'd446,  14'd994,  -14'd259,  -14'd2298,  -14'd35,  14'd184,  14'd1977,  14'd426,  -14'd1181,  
14'd319,  14'd922,  14'd621,  -14'd61,  14'd276,  -14'd1081,  14'd291,  14'd1294,  14'd854,  14'd603,  -14'd1303,  -14'd531,  -14'd1221,  14'd565,  -14'd418,  14'd729,  
14'd291,  14'd1411,  14'd182,  -14'd843,  -14'd742,  14'd787,  -14'd1528,  14'd744,  -14'd711,  -14'd350,  -14'd1201,  -14'd1789,  14'd607,  14'd580,  14'd388,  -14'd234,  
14'd620,  14'd2013,  -14'd39,  -14'd168,  14'd1485,  14'd203,  14'd255,  14'd28,  -14'd1202,  14'd1085,  14'd1388,  -14'd66,  14'd434,  14'd983,  14'd883,  14'd229,  
14'd1109,  -14'd652,  14'd1267,  14'd1196,  14'd1203,  14'd1166,  14'd711,  14'd1482,  -14'd786,  -14'd993,  14'd438,  -14'd720,  14'd257,  -14'd593,  14'd464,  14'd584,  
-14'd1949,  -14'd278,  14'd695,  14'd1170,  14'd272,  14'd1409,  14'd18,  14'd634,  -14'd2072,  -14'd461,  -14'd573,  -14'd537,  -14'd319,  14'd997,  -14'd811,  -14'd911,  
-14'd1083,  14'd418,  14'd565,  14'd653,  14'd437,  -14'd642,  -14'd1541,  14'd483,  -14'd3839,  14'd76,  14'd820,  -14'd420,  14'd67,  -14'd477,  -14'd330,  -14'd1656,  
14'd225,  14'd622,  14'd237,  14'd422,  -14'd1156,  -14'd129,  14'd34,  -14'd52,  -14'd2259,  -14'd370,  14'd1136,  14'd381,  -14'd1356,  -14'd1534,  14'd485,  -14'd905,  
-14'd437,  14'd142,  -14'd641,  -14'd372,  -14'd1077,  14'd913,  14'd897,  14'd644,  14'd492,  -14'd1704,  14'd1221,  14'd1243,  14'd574,  -14'd621,  -14'd293,  14'd171,  
-14'd447,  -14'd382,  14'd258,  -14'd503,  -14'd346,  14'd565,  14'd1442,  14'd1304,  14'd19,  -14'd2198,  -14'd513,  -14'd1298,  -14'd367,  14'd133,  -14'd742,  -14'd170,  
-14'd920,  14'd1410,  -14'd387,  14'd968,  14'd1362,  14'd692,  -14'd1374,  14'd426,  14'd578,  14'd43,  14'd1148,  -14'd154,  14'd77,  -14'd1429,  -14'd195,  -14'd138,  
-14'd1344,  14'd1020,  -14'd394,  14'd1386,  14'd976,  14'd162,  14'd1048,  14'd657,  14'd1638,  -14'd542,  14'd707,  -14'd9,  -14'd843,  -14'd1550,  14'd39,  -14'd346,  
14'd723,  14'd46,  -14'd519,  14'd1369,  14'd786,  -14'd818,  14'd1652,  14'd511,  14'd1720,  -14'd64,  -14'd341,  14'd81,  -14'd140,  -14'd162,  -14'd692,  -14'd723,  
14'd156,  -14'd73,  -14'd125,  14'd237,  -14'd156,  -14'd517,  -14'd584,  14'd618,  14'd676,  14'd1196,  -14'd1260,  14'd87,  14'd990,  14'd1053,  14'd379,  -14'd968,  
-14'd462,  14'd96,  -14'd1448,  -14'd2488,  -14'd947,  14'd334,  -14'd1295,  -14'd1455,  -14'd394,  -14'd785,  14'd332,  -14'd490,  -14'd884,  14'd810,  -14'd1547,  -14'd233,  

-14'd103,  14'd1095,  -14'd1570,  -14'd647,  -14'd1121,  14'd368,  -14'd320,  -14'd163,  -14'd324,  14'd66,  14'd1073,  -14'd802,  -14'd985,  -14'd342,  14'd151,  14'd366,  
14'd274,  14'd337,  -14'd247,  14'd93,  -14'd862,  14'd1649,  14'd932,  -14'd932,  -14'd267,  -14'd1351,  -14'd408,  14'd168,  -14'd1167,  14'd147,  -14'd1814,  14'd591,  
-14'd1212,  -14'd1289,  -14'd1250,  -14'd962,  14'd861,  14'd251,  14'd538,  14'd731,  14'd527,  14'd912,  14'd459,  14'd1203,  14'd35,  14'd387,  14'd1287,  -14'd788,  
14'd372,  14'd451,  14'd869,  -14'd1192,  -14'd688,  -14'd977,  -14'd338,  14'd656,  14'd1254,  14'd678,  -14'd56,  -14'd37,  -14'd463,  14'd1544,  -14'd451,  14'd654,  
-14'd368,  14'd1101,  14'd335,  14'd787,  14'd746,  14'd206,  14'd1287,  -14'd582,  14'd725,  14'd1178,  14'd860,  14'd826,  -14'd586,  -14'd465,  -14'd18,  -14'd1512,  
14'd580,  -14'd172,  14'd275,  14'd701,  -14'd927,  14'd190,  14'd883,  -14'd90,  14'd1471,  14'd1808,  -14'd282,  14'd776,  -14'd377,  -14'd93,  -14'd703,  -14'd1248,  
14'd168,  14'd516,  14'd555,  -14'd915,  14'd57,  14'd903,  14'd1692,  14'd192,  14'd1054,  -14'd942,  -14'd101,  14'd490,  -14'd423,  14'd1647,  -14'd160,  14'd1093,  
-14'd118,  -14'd57,  14'd1406,  -14'd1009,  -14'd817,  -14'd721,  14'd21,  -14'd84,  14'd187,  14'd762,  14'd287,  -14'd342,  -14'd257,  14'd231,  14'd540,  -14'd830,  
14'd1121,  14'd737,  14'd463,  14'd322,  -14'd344,  -14'd781,  -14'd1408,  -14'd1953,  -14'd210,  -14'd42,  -14'd802,  -14'd321,  -14'd1305,  14'd1155,  14'd338,  14'd234,  
-14'd42,  -14'd394,  -14'd1356,  -14'd134,  -14'd1476,  14'd1231,  14'd3,  -14'd184,  14'd1120,  -14'd1040,  14'd667,  -14'd199,  14'd346,  14'd299,  14'd660,  -14'd874,  
14'd1101,  -14'd546,  14'd584,  14'd832,  14'd542,  -14'd299,  14'd293,  -14'd6,  14'd215,  -14'd910,  -14'd1407,  14'd619,  14'd1977,  14'd496,  14'd141,  14'd725,  
14'd363,  14'd1408,  14'd42,  14'd23,  14'd1301,  14'd15,  14'd297,  14'd659,  -14'd109,  14'd394,  14'd1516,  14'd1280,  -14'd121,  14'd1688,  -14'd465,  -14'd433,  
-14'd43,  14'd537,  -14'd282,  -14'd168,  -14'd334,  14'd763,  14'd24,  14'd1030,  -14'd1776,  -14'd824,  -14'd111,  14'd590,  -14'd240,  14'd358,  -14'd140,  -14'd404,  
14'd2279,  14'd961,  14'd103,  14'd896,  -14'd168,  -14'd294,  14'd484,  14'd673,  -14'd996,  -14'd2266,  -14'd148,  -14'd102,  14'd66,  14'd672,  14'd939,  -14'd1155,  
14'd349,  -14'd12,  -14'd1814,  -14'd1103,  -14'd750,  14'd398,  -14'd275,  -14'd386,  14'd1036,  -14'd1018,  -14'd608,  -14'd614,  14'd1003,  14'd481,  -14'd98,  14'd1494,  
14'd179,  14'd808,  -14'd85,  -14'd619,  14'd1779,  14'd545,  -14'd271,  14'd503,  -14'd1285,  -14'd287,  14'd273,  -14'd41,  -14'd20,  14'd1259,  -14'd11,  14'd1260,  
-14'd338,  -14'd740,  -14'd640,  -14'd376,  14'd2164,  -14'd1699,  -14'd294,  14'd333,  -14'd361,  -14'd414,  -14'd175,  -14'd182,  14'd1082,  -14'd764,  -14'd777,  -14'd57,  
14'd678,  14'd1241,  -14'd1326,  14'd17,  14'd108,  -14'd88,  14'd633,  -14'd407,  14'd995,  -14'd36,  -14'd1694,  14'd173,  -14'd1056,  14'd806,  -14'd1173,  14'd1193,  
14'd161,  -14'd301,  14'd206,  -14'd488,  -14'd641,  14'd459,  -14'd939,  14'd710,  -14'd756,  -14'd243,  -14'd1175,  -14'd118,  14'd1173,  14'd265,  -14'd1053,  -14'd261,  
14'd3,  -14'd1368,  -14'd681,  -14'd433,  -14'd968,  -14'd933,  14'd1256,  -14'd1178,  -14'd416,  -14'd1708,  14'd514,  14'd939,  14'd1124,  -14'd193,  14'd17,  14'd608,  
14'd441,  14'd1280,  14'd1432,  14'd215,  -14'd1037,  14'd399,  -14'd1453,  14'd815,  -14'd2461,  -14'd190,  14'd729,  -14'd22,  14'd588,  -14'd979,  -14'd335,  -14'd212,  
-14'd1309,  -14'd851,  14'd64,  -14'd1338,  14'd948,  -14'd1233,  14'd962,  14'd773,  14'd1100,  -14'd1785,  -14'd1419,  14'd105,  14'd662,  14'd850,  -14'd1535,  -14'd389,  
-14'd2069,  -14'd361,  -14'd933,  -14'd817,  -14'd192,  14'd641,  -14'd348,  14'd840,  14'd660,  -14'd1357,  -14'd578,  -14'd815,  -14'd412,  14'd1841,  14'd314,  14'd350,  
-14'd1278,  -14'd1242,  14'd1146,  -14'd224,  14'd376,  -14'd1132,  14'd735,  -14'd328,  -14'd529,  -14'd402,  -14'd1677,  -14'd750,  14'd177,  14'd1466,  -14'd1115,  14'd35,  
14'd44,  -14'd315,  -14'd1498,  14'd83,  14'd396,  -14'd25,  14'd3,  14'd1103,  -14'd1866,  -14'd98,  -14'd956,  14'd297,  14'd692,  -14'd982,  14'd134,  -14'd477,  

14'd613,  14'd822,  14'd561,  14'd146,  -14'd807,  14'd137,  -14'd1689,  -14'd9,  14'd753,  -14'd927,  -14'd1226,  14'd1102,  14'd872,  -14'd383,  -14'd807,  14'd761,  
14'd58,  -14'd182,  -14'd237,  14'd932,  -14'd184,  -14'd403,  -14'd1218,  -14'd189,  -14'd203,  14'd737,  14'd1047,  14'd299,  14'd1012,  14'd2437,  -14'd1443,  -14'd1594,  
-14'd1232,  14'd1215,  14'd534,  -14'd786,  -14'd865,  14'd30,  -14'd1272,  -14'd924,  14'd1389,  -14'd498,  -14'd653,  -14'd260,  -14'd812,  14'd1171,  14'd581,  -14'd158,  
14'd56,  14'd242,  -14'd248,  14'd409,  -14'd926,  14'd280,  -14'd1180,  14'd249,  -14'd493,  -14'd524,  -14'd1345,  14'd59,  -14'd937,  14'd767,  14'd1707,  14'd756,  
14'd1320,  14'd382,  -14'd1570,  14'd1707,  14'd709,  -14'd523,  -14'd397,  14'd438,  14'd1112,  14'd692,  14'd525,  14'd188,  14'd1157,  14'd1223,  14'd1131,  14'd503,  
14'd838,  -14'd1263,  14'd544,  14'd813,  -14'd1709,  14'd1191,  -14'd783,  14'd1362,  -14'd230,  14'd250,  -14'd1487,  14'd160,  -14'd96,  14'd692,  14'd320,  14'd192,  
-14'd485,  -14'd2179,  14'd1646,  -14'd454,  14'd458,  14'd623,  14'd968,  -14'd322,  -14'd519,  -14'd636,  14'd537,  -14'd906,  14'd15,  14'd962,  14'd1409,  14'd445,  
14'd753,  -14'd79,  -14'd128,  -14'd189,  -14'd988,  14'd491,  14'd378,  -14'd1241,  -14'd419,  14'd1151,  -14'd1090,  -14'd313,  -14'd1235,  14'd1881,  14'd658,  -14'd1433,  
-14'd272,  14'd550,  -14'd175,  -14'd171,  14'd79,  -14'd730,  14'd85,  -14'd283,  14'd1120,  -14'd406,  14'd282,  14'd1128,  -14'd811,  -14'd1389,  14'd5,  -14'd482,  
14'd840,  14'd1126,  -14'd490,  -14'd435,  -14'd1609,  14'd1453,  -14'd502,  -14'd697,  14'd1803,  14'd32,  14'd821,  14'd212,  14'd294,  14'd1712,  -14'd1069,  14'd1897,  
-14'd60,  14'd244,  -14'd12,  14'd1633,  -14'd956,  14'd615,  14'd38,  14'd815,  14'd306,  14'd952,  14'd1467,  -14'd397,  14'd274,  -14'd679,  14'd262,  -14'd196,  
14'd330,  14'd1224,  14'd3,  14'd599,  14'd686,  14'd487,  -14'd87,  14'd1152,  -14'd442,  14'd1152,  -14'd811,  -14'd526,  -14'd583,  14'd1324,  -14'd94,  14'd998,  
-14'd1206,  14'd64,  -14'd240,  -14'd1603,  14'd1289,  14'd608,  14'd737,  14'd26,  -14'd856,  -14'd271,  14'd706,  -14'd611,  -14'd604,  14'd440,  -14'd666,  14'd117,  
-14'd1773,  14'd1249,  -14'd348,  -14'd646,  14'd834,  -14'd1026,  -14'd532,  -14'd230,  -14'd1128,  -14'd115,  -14'd670,  14'd1601,  -14'd1815,  -14'd452,  14'd1087,  14'd871,  
-14'd794,  14'd900,  14'd678,  14'd804,  14'd225,  14'd580,  14'd271,  14'd851,  14'd509,  -14'd153,  -14'd736,  -14'd498,  -14'd1349,  -14'd44,  -14'd477,  -14'd158,  
-14'd474,  14'd1087,  14'd1042,  14'd109,  14'd76,  14'd739,  14'd723,  14'd1345,  14'd301,  -14'd565,  -14'd22,  14'd648,  14'd961,  -14'd1424,  14'd506,  -14'd128,  
14'd608,  14'd320,  14'd338,  -14'd808,  14'd1520,  -14'd791,  -14'd357,  -14'd328,  -14'd532,  14'd824,  14'd52,  14'd276,  14'd288,  14'd130,  14'd1399,  -14'd591,  
14'd432,  -14'd193,  -14'd820,  -14'd104,  14'd253,  14'd98,  -14'd949,  14'd493,  -14'd1778,  -14'd991,  14'd1679,  14'd270,  14'd795,  14'd1175,  -14'd1040,  -14'd285,  
14'd363,  14'd1002,  14'd507,  14'd1150,  14'd960,  14'd581,  14'd30,  14'd1646,  14'd630,  -14'd483,  -14'd193,  14'd981,  14'd444,  14'd538,  -14'd98,  -14'd91,  
14'd2007,  14'd226,  -14'd406,  14'd753,  -14'd691,  -14'd104,  -14'd1345,  14'd727,  14'd947,  14'd485,  -14'd4,  -14'd414,  -14'd785,  14'd812,  14'd298,  -14'd267,  
-14'd1310,  14'd542,  -14'd1235,  -14'd704,  -14'd1400,  14'd912,  14'd2084,  14'd84,  14'd1260,  -14'd753,  14'd34,  -14'd442,  -14'd1140,  -14'd307,  -14'd65,  14'd1098,  
-14'd1025,  -14'd632,  -14'd375,  -14'd991,  14'd699,  14'd1501,  14'd424,  14'd423,  14'd267,  14'd96,  14'd1150,  14'd71,  14'd1093,  -14'd1324,  14'd1684,  -14'd346,  
14'd971,  -14'd318,  -14'd1906,  -14'd1670,  14'd530,  -14'd79,  -14'd508,  14'd94,  14'd115,  14'd509,  14'd227,  14'd1020,  14'd137,  14'd304,  -14'd1259,  -14'd1088,  
14'd2268,  14'd1881,  14'd143,  14'd414,  14'd1208,  14'd116,  14'd69,  14'd158,  -14'd405,  14'd1499,  14'd619,  14'd712,  -14'd22,  14'd1218,  14'd1246,  -14'd176,  
-14'd895,  14'd1571,  -14'd569,  14'd985,  -14'd548,  14'd398,  14'd963,  14'd1957,  14'd874,  -14'd1437,  -14'd813,  14'd1768,  -14'd304,  -14'd953,  14'd626,  14'd1115,  

-14'd544,  14'd945,  -14'd731,  -14'd272,  14'd1138,  14'd755,  -14'd267,  14'd440,  14'd488,  -14'd37,  -14'd1442,  -14'd274,  14'd348,  14'd565,  -14'd1196,  14'd1262,  
14'd824,  14'd803,  -14'd1234,  -14'd701,  14'd229,  14'd567,  14'd97,  14'd705,  -14'd1610,  -14'd725,  -14'd835,  -14'd890,  14'd317,  14'd206,  -14'd817,  -14'd944,  
-14'd989,  14'd863,  -14'd252,  14'd1160,  -14'd774,  -14'd116,  14'd476,  -14'd90,  14'd334,  -14'd56,  -14'd50,  -14'd368,  14'd133,  14'd1248,  14'd922,  -14'd1249,  
14'd1048,  -14'd89,  -14'd1104,  -14'd678,  -14'd457,  14'd233,  14'd768,  -14'd1056,  14'd78,  14'd683,  14'd620,  -14'd1451,  -14'd704,  14'd316,  14'd56,  -14'd79,  
14'd611,  -14'd749,  14'd1385,  14'd344,  14'd752,  -14'd1046,  -14'd398,  14'd214,  -14'd1204,  14'd265,  -14'd1024,  -14'd523,  -14'd78,  -14'd1251,  -14'd295,  14'd956,  
14'd131,  -14'd459,  14'd1010,  -14'd24,  -14'd579,  -14'd282,  14'd654,  -14'd796,  -14'd59,  -14'd507,  14'd71,  14'd206,  -14'd613,  -14'd453,  14'd520,  -14'd156,  
-14'd349,  -14'd53,  -14'd953,  14'd603,  14'd277,  -14'd47,  -14'd330,  -14'd345,  -14'd690,  14'd461,  14'd373,  14'd898,  -14'd1090,  14'd1308,  -14'd242,  -14'd624,  
14'd125,  -14'd387,  14'd94,  -14'd1760,  14'd550,  -14'd28,  14'd157,  -14'd1543,  14'd383,  -14'd29,  -14'd620,  14'd280,  -14'd1144,  14'd480,  14'd284,  -14'd705,  
-14'd86,  -14'd90,  14'd515,  14'd177,  14'd163,  -14'd1386,  -14'd567,  -14'd671,  -14'd28,  -14'd673,  14'd309,  14'd254,  -14'd30,  14'd476,  14'd170,  14'd109,  
14'd370,  -14'd831,  14'd526,  14'd613,  14'd435,  14'd359,  -14'd584,  14'd298,  14'd1421,  14'd351,  14'd243,  14'd64,  -14'd103,  14'd849,  -14'd527,  -14'd1069,  
-14'd208,  -14'd869,  -14'd622,  14'd150,  -14'd473,  14'd514,  14'd662,  -14'd1699,  -14'd180,  14'd529,  -14'd285,  14'd13,  14'd561,  14'd692,  14'd1080,  -14'd1168,  
14'd27,  -14'd87,  -14'd1290,  -14'd336,  -14'd858,  -14'd1042,  14'd980,  -14'd877,  -14'd1561,  -14'd190,  14'd259,  -14'd442,  -14'd626,  14'd57,  -14'd1442,  -14'd492,  
-14'd340,  14'd945,  14'd901,  14'd48,  -14'd624,  -14'd299,  -14'd790,  14'd424,  -14'd1095,  -14'd1586,  -14'd200,  14'd499,  14'd322,  14'd307,  -14'd1231,  14'd797,  
-14'd309,  -14'd1395,  14'd22,  -14'd472,  14'd178,  -14'd60,  14'd1046,  -14'd1069,  -14'd785,  -14'd493,  -14'd1416,  14'd196,  -14'd648,  14'd1079,  -14'd1150,  -14'd1009,  
-14'd604,  -14'd1480,  -14'd539,  14'd3,  -14'd775,  14'd696,  -14'd654,  14'd335,  -14'd211,  -14'd1061,  14'd264,  -14'd1360,  -14'd917,  -14'd507,  14'd1127,  14'd185,  
-14'd88,  14'd601,  14'd1203,  -14'd1131,  -14'd400,  14'd1143,  -14'd1543,  -14'd106,  -14'd1283,  -14'd1115,  14'd686,  -14'd1271,  14'd291,  14'd1298,  14'd687,  -14'd215,  
-14'd1079,  -14'd894,  14'd236,  -14'd933,  -14'd1035,  14'd31,  14'd1367,  -14'd467,  14'd497,  14'd557,  14'd287,  14'd249,  -14'd202,  14'd1161,  -14'd334,  14'd152,  
-14'd327,  14'd479,  -14'd1035,  -14'd1077,  14'd189,  -14'd121,  -14'd1115,  14'd207,  -14'd340,  -14'd27,  14'd666,  14'd842,  -14'd900,  -14'd816,  -14'd1034,  -14'd431,  
-14'd1467,  -14'd380,  -14'd847,  14'd459,  14'd208,  14'd963,  -14'd125,  -14'd101,  -14'd353,  14'd365,  14'd594,  -14'd271,  -14'd219,  14'd176,  -14'd194,  -14'd797,  
-14'd828,  -14'd1126,  14'd482,  14'd106,  14'd800,  14'd267,  14'd154,  -14'd194,  14'd403,  -14'd505,  -14'd1386,  14'd627,  -14'd497,  14'd84,  -14'd737,  14'd414,  
-14'd111,  -14'd335,  14'd517,  14'd1440,  14'd471,  -14'd806,  14'd454,  14'd21,  -14'd109,  14'd850,  14'd118,  -14'd26,  14'd199,  -14'd883,  -14'd867,  -14'd483,  
-14'd951,  -14'd138,  14'd1269,  -14'd227,  -14'd353,  -14'd44,  -14'd992,  14'd65,  -14'd820,  14'd209,  14'd1011,  -14'd169,  14'd213,  -14'd64,  -14'd322,  14'd654,  
-14'd375,  -14'd222,  14'd76,  -14'd337,  14'd466,  14'd762,  -14'd972,  14'd121,  14'd629,  -14'd885,  -14'd749,  -14'd1284,  -14'd498,  -14'd1499,  -14'd1386,  -14'd198,  
-14'd328,  14'd1359,  -14'd770,  14'd128,  -14'd351,  -14'd502,  14'd12,  14'd86,  14'd623,  14'd736,  -14'd910,  -14'd547,  -14'd1698,  -14'd319,  -14'd760,  -14'd1614,  
-14'd1221,  14'd314,  -14'd470,  -14'd424,  -14'd1360,  14'd571,  -14'd1129,  14'd859,  -14'd632,  14'd1070,  -14'd490,  -14'd924,  14'd26,  -14'd373,  -14'd1536,  14'd213,  

-14'd560,  -14'd249,  14'd1142,  -14'd1074,  -14'd940,  14'd903,  14'd4,  -14'd1135,  -14'd598,  14'd258,  14'd452,  -14'd406,  14'd151,  14'd1113,  -14'd1067,  -14'd769,  
-14'd187,  14'd182,  14'd886,  14'd512,  -14'd416,  -14'd69,  14'd686,  14'd535,  14'd570,  -14'd794,  -14'd75,  14'd1270,  14'd508,  14'd1076,  -14'd384,  -14'd179,  
14'd1072,  14'd328,  14'd632,  14'd442,  14'd97,  14'd235,  14'd613,  -14'd79,  14'd275,  -14'd778,  -14'd264,  -14'd746,  14'd1214,  -14'd256,  -14'd648,  14'd246,  
14'd1456,  -14'd161,  -14'd1266,  -14'd74,  -14'd935,  14'd294,  14'd1262,  14'd539,  -14'd242,  -14'd1290,  14'd152,  -14'd281,  14'd790,  -14'd2467,  -14'd840,  14'd1246,  
14'd1032,  14'd1706,  -14'd749,  14'd1149,  14'd95,  -14'd311,  14'd1223,  -14'd423,  14'd461,  14'd347,  -14'd48,  14'd1068,  14'd1135,  14'd1352,  14'd228,  14'd2456,  
14'd386,  14'd315,  14'd780,  -14'd117,  -14'd718,  14'd949,  -14'd289,  -14'd655,  -14'd324,  14'd349,  -14'd539,  14'd1421,  14'd692,  14'd371,  -14'd648,  14'd1413,  
-14'd646,  14'd692,  14'd626,  14'd1147,  -14'd1330,  14'd665,  14'd305,  14'd595,  14'd983,  -14'd1447,  -14'd260,  14'd201,  -14'd829,  -14'd905,  -14'd507,  -14'd284,  
-14'd803,  14'd496,  -14'd728,  14'd150,  14'd1392,  -14'd10,  -14'd520,  14'd1337,  -14'd24,  14'd317,  -14'd951,  -14'd131,  14'd1535,  -14'd528,  -14'd1504,  -14'd340,  
14'd269,  14'd371,  -14'd1612,  14'd691,  14'd671,  -14'd462,  -14'd1489,  14'd397,  14'd335,  14'd1518,  14'd1480,  -14'd307,  14'd574,  -14'd2196,  14'd1470,  14'd972,  
-14'd203,  -14'd2149,  -14'd787,  14'd1849,  14'd1607,  14'd946,  -14'd474,  -14'd434,  14'd90,  -14'd596,  14'd774,  14'd170,  14'd926,  14'd652,  14'd621,  14'd1031,  
-14'd858,  14'd306,  -14'd328,  -14'd522,  -14'd1780,  -14'd1445,  14'd1301,  14'd487,  14'd345,  14'd232,  -14'd1992,  14'd193,  -14'd733,  14'd239,  14'd1880,  14'd834,  
-14'd1319,  14'd439,  -14'd422,  -14'd573,  -14'd212,  -14'd123,  14'd463,  14'd969,  14'd34,  14'd256,  -14'd723,  -14'd187,  -14'd1792,  -14'd170,  14'd881,  -14'd1126,  
-14'd911,  -14'd260,  14'd1680,  14'd1667,  -14'd1004,  -14'd723,  14'd14,  -14'd71,  14'd721,  14'd1451,  -14'd1252,  -14'd723,  -14'd647,  14'd425,  14'd1053,  -14'd264,  
-14'd450,  14'd358,  -14'd2097,  -14'd430,  14'd1063,  14'd307,  14'd895,  14'd270,  -14'd761,  14'd98,  -14'd386,  -14'd669,  14'd1726,  -14'd1270,  14'd933,  14'd1324,  
-14'd2473,  -14'd995,  14'd14,  -14'd328,  14'd1034,  -14'd1292,  -14'd1196,  -14'd119,  14'd1078,  14'd298,  14'd695,  -14'd773,  -14'd1761,  -14'd608,  -14'd75,  14'd1154,  
-14'd911,  14'd1088,  14'd322,  14'd1372,  -14'd368,  -14'd591,  -14'd496,  -14'd180,  -14'd661,  14'd139,  -14'd2735,  -14'd167,  14'd208,  -14'd103,  14'd638,  14'd259,  
-14'd572,  -14'd1005,  14'd708,  14'd35,  14'd671,  14'd1127,  14'd54,  -14'd348,  -14'd2297,  14'd660,  -14'd1552,  -14'd834,  14'd1512,  14'd40,  14'd455,  -14'd599,  
-14'd1048,  14'd664,  14'd734,  -14'd478,  14'd1053,  -14'd155,  -14'd769,  -14'd568,  -14'd1033,  14'd587,  14'd1363,  14'd1507,  14'd356,  14'd1920,  -14'd1349,  14'd515,  
-14'd662,  -14'd759,  14'd921,  14'd583,  14'd450,  -14'd166,  14'd730,  -14'd966,  -14'd310,  -14'd210,  14'd2076,  -14'd718,  -14'd254,  -14'd855,  14'd235,  14'd458,  
14'd152,  14'd1282,  14'd110,  -14'd384,  14'd927,  14'd546,  14'd561,  14'd32,  14'd677,  -14'd584,  -14'd616,  14'd530,  -14'd40,  14'd466,  14'd162,  14'd142,  
-14'd585,  14'd820,  -14'd1813,  -14'd74,  -14'd676,  -14'd317,  14'd541,  14'd296,  14'd1250,  14'd422,  -14'd1342,  -14'd212,  -14'd322,  14'd50,  -14'd675,  -14'd1090,  
14'd587,  14'd716,  14'd621,  -14'd369,  -14'd93,  -14'd602,  14'd568,  14'd406,  14'd62,  -14'd1139,  -14'd795,  14'd1849,  -14'd675,  -14'd302,  14'd592,  14'd278,  
-14'd1410,  14'd954,  -14'd1320,  -14'd473,  -14'd1227,  -14'd982,  14'd1480,  -14'd78,  14'd285,  14'd744,  -14'd447,  -14'd451,  14'd581,  14'd469,  14'd505,  -14'd19,  
14'd407,  -14'd38,  14'd67,  -14'd555,  -14'd698,  -14'd1129,  14'd180,  14'd916,  14'd647,  -14'd1023,  14'd963,  14'd396,  -14'd1206,  14'd1217,  -14'd198,  -14'd413,  
14'd1397,  -14'd597,  -14'd1615,  -14'd493,  14'd37,  14'd314,  14'd1468,  14'd751,  -14'd637,  -14'd1525,  -14'd16,  -14'd810,  -14'd825,  14'd1964,  -14'd147,  -14'd1484,  

-14'd1277,  -14'd965,  -14'd1668,  -14'd545,  -14'd443,  -14'd687,  14'd2721,  -14'd1318,  14'd154,  14'd943,  -14'd383,  -14'd945,  -14'd568,  -14'd836,  -14'd1242,  -14'd1099,  
14'd312,  -14'd1117,  14'd164,  14'd155,  -14'd474,  14'd12,  14'd236,  14'd244,  14'd1464,  14'd672,  -14'd259,  -14'd680,  -14'd474,  14'd802,  -14'd1748,  14'd61,  
14'd880,  14'd278,  -14'd883,  -14'd1653,  14'd367,  -14'd153,  -14'd952,  -14'd805,  14'd351,  -14'd869,  14'd452,  -14'd1313,  14'd732,  -14'd455,  -14'd35,  14'd751,  
14'd932,  14'd1092,  14'd464,  14'd645,  14'd888,  14'd420,  -14'd963,  -14'd107,  14'd411,  14'd1240,  14'd136,  14'd242,  -14'd526,  -14'd412,  14'd1397,  -14'd52,  
-14'd2029,  -14'd346,  14'd1541,  14'd391,  14'd233,  14'd107,  -14'd188,  -14'd67,  -14'd1112,  14'd1527,  -14'd9,  -14'd72,  -14'd123,  -14'd523,  14'd580,  -14'd707,  
-14'd815,  14'd98,  14'd1343,  14'd359,  -14'd1066,  14'd422,  14'd288,  -14'd486,  -14'd470,  -14'd723,  14'd204,  -14'd221,  -14'd1187,  -14'd899,  -14'd60,  -14'd226,  
14'd879,  14'd562,  -14'd586,  14'd1759,  -14'd1456,  14'd1461,  -14'd1288,  -14'd1724,  14'd880,  -14'd170,  14'd433,  -14'd465,  14'd31,  -14'd1443,  -14'd1523,  -14'd397,  
-14'd36,  -14'd364,  14'd168,  14'd353,  14'd549,  -14'd560,  14'd288,  -14'd1155,  -14'd202,  -14'd592,  14'd1405,  -14'd415,  14'd875,  -14'd720,  -14'd956,  14'd1626,  
-14'd1154,  14'd1038,  14'd389,  14'd640,  14'd567,  -14'd670,  14'd199,  14'd376,  -14'd316,  14'd414,  14'd173,  -14'd1195,  -14'd461,  14'd841,  -14'd612,  14'd392,  
-14'd102,  -14'd318,  14'd1606,  14'd515,  14'd435,  14'd1182,  -14'd559,  14'd547,  -14'd385,  14'd646,  -14'd1416,  14'd1241,  -14'd830,  14'd405,  -14'd180,  -14'd1563,  
14'd788,  14'd1143,  -14'd768,  14'd1195,  -14'd2969,  -14'd1345,  14'd676,  14'd94,  14'd15,  14'd206,  -14'd1637,  14'd469,  14'd77,  -14'd823,  -14'd227,  -14'd36,  
14'd509,  14'd320,  14'd583,  -14'd259,  -14'd1021,  -14'd427,  14'd683,  14'd519,  14'd2474,  -14'd860,  14'd919,  -14'd915,  14'd187,  14'd1145,  -14'd395,  14'd660,  
-14'd1091,  14'd794,  -14'd163,  14'd788,  14'd1826,  -14'd581,  14'd1009,  14'd243,  14'd532,  14'd99,  14'd26,  14'd277,  14'd166,  -14'd107,  -14'd1189,  -14'd614,  
14'd1345,  -14'd426,  -14'd514,  -14'd319,  14'd522,  -14'd1043,  -14'd403,  14'd1044,  -14'd1782,  -14'd181,  14'd515,  14'd737,  -14'd789,  14'd789,  14'd1307,  -14'd1169,  
14'd205,  14'd282,  14'd1308,  14'd469,  14'd311,  14'd312,  -14'd365,  14'd647,  14'd1560,  14'd367,  14'd276,  14'd205,  14'd1312,  14'd772,  14'd1156,  14'd460,  
-14'd68,  -14'd542,  14'd774,  14'd37,  -14'd958,  -14'd126,  14'd766,  14'd517,  14'd200,  -14'd366,  -14'd286,  14'd675,  14'd226,  14'd1238,  14'd1289,  -14'd956,  
14'd217,  14'd462,  14'd423,  14'd977,  -14'd811,  14'd240,  14'd396,  14'd79,  14'd1088,  -14'd885,  14'd1053,  -14'd191,  -14'd943,  -14'd520,  -14'd653,  -14'd1086,  
-14'd1042,  -14'd1299,  -14'd1131,  -14'd710,  -14'd40,  14'd1350,  14'd834,  -14'd1320,  -14'd210,  14'd723,  14'd1794,  -14'd560,  -14'd491,  -14'd971,  -14'd321,  14'd827,  
-14'd973,  14'd1180,  -14'd766,  -14'd942,  14'd82,  14'd1127,  14'd257,  -14'd189,  -14'd506,  14'd1355,  14'd270,  -14'd429,  14'd1532,  14'd264,  -14'd303,  14'd22,  
14'd267,  -14'd382,  14'd352,  14'd78,  14'd952,  14'd1283,  -14'd1234,  14'd807,  14'd316,  14'd812,  14'd136,  14'd565,  14'd847,  -14'd1203,  14'd1175,  14'd2221,  
-14'd451,  -14'd1352,  14'd1198,  14'd374,  14'd1018,  -14'd341,  -14'd1732,  14'd1168,  -14'd29,  -14'd633,  14'd41,  -14'd24,  -14'd433,  14'd1608,  14'd1506,  -14'd193,  
-14'd1926,  -14'd901,  -14'd231,  14'd577,  14'd32,  14'd710,  -14'd201,  14'd1174,  -14'd609,  -14'd731,  14'd409,  -14'd105,  14'd519,  -14'd797,  14'd19,  -14'd1018,  
-14'd752,  -14'd2850,  -14'd602,  14'd476,  14'd272,  14'd768,  -14'd1123,  -14'd839,  -14'd1277,  -14'd156,  14'd752,  -14'd809,  14'd151,  -14'd1229,  -14'd261,  14'd1253,  
-14'd431,  14'd256,  14'd245,  -14'd1237,  14'd903,  -14'd1036,  14'd251,  14'd190,  14'd150,  14'd1795,  14'd580,  14'd348,  -14'd504,  -14'd1231,  14'd507,  -14'd677,  
-14'd1523,  14'd266,  -14'd1258,  -14'd1297,  14'd1016,  -14'd1464,  -14'd925,  -14'd434,  14'd1297,  14'd2261,  -14'd342,  14'd390,  14'd916,  -14'd2110,  14'd16,  -14'd716,  

-14'd1238,  -14'd964,  14'd277,  -14'd636,  -14'd1430,  14'd286,  -14'd1755,  -14'd451,  -14'd1077,  -14'd531,  -14'd783,  -14'd966,  14'd447,  14'd1417,  14'd645,  14'd227,  
14'd15,  -14'd126,  14'd9,  -14'd908,  14'd1,  14'd214,  -14'd198,  14'd870,  -14'd1079,  14'd1745,  -14'd370,  -14'd578,  14'd1236,  -14'd399,  -14'd1425,  14'd720,  
-14'd645,  -14'd1249,  14'd38,  -14'd889,  14'd150,  14'd1009,  -14'd180,  14'd1152,  14'd480,  -14'd384,  -14'd492,  -14'd33,  14'd1563,  -14'd601,  14'd836,  -14'd613,  
-14'd508,  14'd1751,  14'd158,  14'd450,  14'd142,  -14'd285,  -14'd1589,  -14'd325,  -14'd408,  -14'd971,  14'd836,  -14'd141,  -14'd239,  -14'd2073,  14'd1670,  -14'd1492,  
14'd1717,  -14'd77,  -14'd65,  14'd1997,  -14'd156,  -14'd178,  -14'd22,  -14'd361,  -14'd736,  -14'd245,  14'd1001,  14'd740,  -14'd808,  -14'd510,  14'd1173,  -14'd744,  
-14'd1085,  -14'd672,  14'd137,  -14'd1796,  -14'd656,  14'd655,  14'd276,  -14'd1217,  14'd513,  -14'd757,  -14'd1020,  -14'd269,  14'd46,  -14'd586,  14'd809,  14'd1273,  
14'd1513,  -14'd544,  14'd216,  14'd879,  -14'd554,  -14'd627,  14'd106,  14'd63,  -14'd970,  -14'd136,  -14'd5,  -14'd432,  14'd678,  14'd259,  14'd39,  14'd209,  
14'd2226,  14'd640,  14'd214,  14'd133,  14'd19,  14'd658,  14'd2814,  14'd65,  14'd276,  -14'd901,  -14'd1744,  -14'd851,  -14'd364,  -14'd81,  14'd766,  -14'd1988,  
14'd1173,  14'd1387,  14'd898,  14'd606,  14'd1572,  14'd19,  -14'd143,  -14'd683,  14'd1888,  14'd975,  14'd893,  14'd1535,  -14'd313,  14'd1462,  14'd1497,  -14'd184,  
14'd170,  -14'd940,  -14'd161,  -14'd336,  -14'd787,  14'd542,  14'd685,  14'd855,  14'd1762,  -14'd126,  14'd768,  14'd1686,  -14'd481,  14'd589,  14'd88,  -14'd1056,  
-14'd1718,  -14'd299,  -14'd386,  14'd192,  -14'd2027,  14'd435,  14'd405,  -14'd770,  -14'd1102,  -14'd1526,  -14'd620,  14'd200,  -14'd811,  14'd1729,  14'd875,  -14'd193,  
14'd2195,  14'd456,  -14'd142,  -14'd755,  -14'd1065,  -14'd185,  -14'd71,  -14'd748,  -14'd201,  -14'd406,  -14'd95,  14'd1554,  14'd251,  14'd325,  -14'd1225,  14'd610,  
14'd770,  14'd1628,  14'd750,  -14'd616,  14'd999,  14'd49,  14'd1847,  -14'd91,  14'd435,  14'd196,  -14'd517,  14'd662,  14'd283,  14'd748,  14'd261,  -14'd285,  
14'd893,  14'd941,  14'd552,  -14'd497,  -14'd508,  14'd755,  -14'd300,  14'd54,  -14'd306,  -14'd1622,  14'd1504,  14'd711,  -14'd701,  -14'd205,  14'd1039,  14'd705,  
14'd457,  14'd885,  -14'd301,  -14'd422,  -14'd609,  -14'd112,  -14'd192,  -14'd1,  14'd2045,  -14'd583,  14'd902,  -14'd671,  -14'd177,  14'd1463,  -14'd58,  -14'd1260,  
14'd181,  -14'd487,  -14'd96,  14'd215,  -14'd589,  -14'd705,  14'd1169,  -14'd1033,  -14'd1257,  -14'd565,  -14'd113,  14'd1148,  14'd484,  -14'd105,  14'd460,  -14'd70,  
14'd1702,  14'd1071,  14'd508,  -14'd334,  -14'd610,  -14'd1018,  14'd681,  14'd171,  -14'd1369,  -14'd1301,  -14'd532,  -14'd85,  14'd860,  -14'd275,  -14'd1161,  14'd191,  
14'd837,  14'd441,  -14'd983,  14'd83,  -14'd1320,  -14'd693,  14'd933,  -14'd441,  -14'd1413,  -14'd770,  14'd1557,  -14'd384,  -14'd321,  14'd1410,  -14'd1399,  -14'd941,  
14'd588,  14'd617,  14'd1357,  -14'd193,  -14'd1259,  14'd659,  14'd971,  14'd300,  -14'd456,  -14'd1523,  14'd1368,  -14'd2,  14'd302,  -14'd1091,  14'd95,  14'd548,  
-14'd916,  -14'd736,  -14'd1739,  -14'd1946,  -14'd352,  -14'd1703,  14'd645,  14'd315,  -14'd1629,  -14'd3208,  -14'd222,  -14'd1810,  14'd592,  14'd361,  -14'd2179,  -14'd152,  
-14'd675,  14'd383,  -14'd273,  -14'd276,  -14'd1630,  -14'd73,  -14'd343,  14'd892,  -14'd977,  14'd646,  14'd1073,  14'd763,  -14'd8,  14'd1077,  14'd840,  -14'd129,  
14'd1020,  -14'd493,  14'd1672,  14'd319,  -14'd430,  -14'd305,  14'd706,  -14'd7,  -14'd1169,  14'd548,  -14'd137,  -14'd990,  14'd436,  14'd633,  14'd385,  14'd704,  
-14'd1104,  14'd1127,  14'd233,  -14'd1164,  14'd313,  -14'd2261,  14'd1290,  -14'd302,  -14'd733,  14'd2078,  -14'd622,  -14'd1373,  -14'd207,  14'd1561,  -14'd1014,  -14'd920,  
-14'd1962,  -14'd1948,  14'd125,  -14'd3238,  -14'd833,  -14'd1474,  14'd136,  -14'd109,  14'd26,  -14'd861,  -14'd1288,  -14'd2099,  -14'd1092,  -14'd53,  -14'd1370,  -14'd778,  
14'd214,  -14'd1343,  -14'd1693,  -14'd2317,  -14'd2165,  -14'd1561,  -14'd1228,  -14'd761,  -14'd1302,  -14'd2516,  -14'd846,  -14'd2416,  -14'd2889,  -14'd746,  -14'd1415,  -14'd2489,  

-14'd228,  14'd560,  14'd923,  14'd366,  -14'd765,  -14'd597,  -14'd136,  -14'd444,  14'd673,  -14'd251,  14'd261,  -14'd388,  14'd753,  14'd401,  -14'd555,  14'd1164,  
14'd298,  14'd1702,  14'd2565,  14'd457,  14'd421,  -14'd645,  14'd980,  14'd344,  14'd1125,  -14'd416,  14'd1005,  14'd542,  14'd310,  14'd64,  -14'd675,  -14'd358,  
-14'd516,  14'd180,  14'd1397,  -14'd234,  14'd923,  14'd1515,  14'd1553,  14'd555,  -14'd234,  -14'd2372,  -14'd338,  14'd1082,  -14'd526,  14'd3106,  14'd856,  -14'd50,  
14'd1070,  14'd34,  14'd127,  14'd409,  14'd963,  -14'd742,  -14'd647,  14'd988,  14'd497,  14'd1494,  14'd674,  14'd799,  -14'd1120,  14'd1182,  14'd184,  14'd1107,  
-14'd1633,  -14'd734,  -14'd7,  14'd1093,  -14'd2602,  -14'd425,  -14'd732,  14'd787,  14'd131,  14'd1036,  -14'd944,  14'd763,  -14'd1299,  -14'd1083,  14'd188,  -14'd1003,  
-14'd672,  14'd1776,  14'd1017,  14'd391,  14'd813,  -14'd620,  14'd992,  -14'd142,  -14'd1636,  -14'd1072,  14'd149,  -14'd1230,  -14'd987,  14'd1168,  -14'd473,  -14'd596,  
14'd660,  -14'd399,  14'd307,  -14'd1125,  14'd19,  14'd69,  14'd720,  -14'd1136,  14'd35,  14'd515,  14'd2242,  14'd78,  14'd1092,  14'd1786,  14'd344,  14'd223,  
-14'd676,  -14'd178,  14'd295,  14'd351,  -14'd892,  14'd762,  14'd337,  -14'd1678,  14'd51,  -14'd455,  14'd432,  14'd30,  14'd943,  14'd495,  -14'd501,  14'd1216,  
-14'd514,  14'd2006,  -14'd1079,  14'd545,  14'd2005,  14'd89,  -14'd1378,  -14'd248,  -14'd386,  14'd407,  -14'd2,  14'd510,  -14'd1042,  -14'd976,  14'd319,  -14'd1342,  
14'd890,  -14'd1988,  14'd413,  -14'd55,  14'd561,  -14'd320,  14'd21,  -14'd1058,  -14'd147,  14'd1417,  -14'd155,  14'd28,  -14'd1081,  14'd398,  14'd575,  -14'd670,  
14'd582,  14'd721,  14'd303,  -14'd1756,  -14'd1966,  -14'd1947,  14'd2163,  -14'd1286,  -14'd1815,  -14'd1192,  14'd1476,  14'd731,  -14'd2073,  14'd1250,  14'd598,  14'd522,  
14'd725,  -14'd375,  14'd1381,  -14'd1127,  -14'd912,  14'd252,  14'd1064,  -14'd224,  14'd83,  -14'd300,  -14'd397,  -14'd432,  -14'd1485,  14'd87,  -14'd617,  -14'd588,  
-14'd369,  14'd1352,  -14'd794,  -14'd2218,  14'd977,  -14'd1256,  14'd353,  14'd581,  14'd1324,  -14'd111,  -14'd716,  -14'd374,  -14'd991,  14'd302,  14'd762,  -14'd82,  
-14'd734,  14'd1730,  -14'd351,  14'd683,  -14'd192,  -14'd909,  14'd1150,  14'd564,  -14'd620,  -14'd975,  14'd269,  -14'd475,  -14'd716,  14'd346,  14'd385,  -14'd616,  
-14'd1626,  14'd313,  14'd228,  -14'd949,  -14'd823,  -14'd908,  14'd471,  -14'd409,  14'd117,  -14'd1445,  -14'd1252,  -14'd31,  -14'd1354,  -14'd740,  14'd727,  14'd615,  
14'd5,  -14'd696,  14'd999,  -14'd711,  -14'd785,  14'd908,  14'd449,  14'd663,  -14'd843,  14'd395,  14'd11,  -14'd429,  -14'd697,  14'd1407,  -14'd638,  -14'd496,  
14'd741,  -14'd249,  14'd511,  -14'd2053,  -14'd793,  -14'd0,  -14'd649,  -14'd512,  14'd582,  -14'd359,  -14'd537,  14'd66,  -14'd1917,  14'd306,  -14'd743,  -14'd1130,  
14'd1390,  -14'd776,  14'd1048,  14'd1017,  -14'd775,  14'd553,  14'd310,  14'd1503,  -14'd1780,  -14'd257,  14'd790,  14'd972,  14'd416,  14'd1668,  14'd1330,  -14'd893,  
-14'd989,  14'd223,  -14'd1194,  14'd2003,  -14'd1179,  -14'd3,  -14'd1077,  -14'd44,  14'd164,  14'd245,  -14'd1416,  -14'd815,  14'd35,  -14'd555,  14'd701,  -14'd980,  
14'd1458,  -14'd55,  14'd1284,  -14'd128,  14'd85,  14'd313,  14'd552,  -14'd538,  14'd749,  14'd965,  14'd32,  14'd1471,  14'd503,  -14'd1030,  -14'd349,  14'd674,  
14'd47,  -14'd1555,  14'd1723,  -14'd1002,  -14'd1561,  -14'd1324,  -14'd1426,  -14'd606,  -14'd1184,  14'd1639,  -14'd2481,  14'd1879,  -14'd136,  14'd1343,  14'd651,  -14'd798,  
14'd189,  14'd1312,  14'd1571,  -14'd921,  -14'd586,  14'd32,  -14'd1145,  14'd1595,  14'd1086,  14'd770,  -14'd1386,  14'd754,  14'd247,  14'd281,  14'd404,  14'd290,  
14'd535,  14'd691,  14'd47,  14'd1832,  14'd593,  14'd2374,  -14'd724,  14'd2063,  14'd1080,  -14'd1932,  -14'd701,  -14'd2062,  14'd1121,  -14'd1032,  14'd98,  14'd336,  
-14'd878,  -14'd962,  14'd713,  -14'd912,  14'd725,  -14'd580,  -14'd1183,  -14'd156,  -14'd1515,  14'd758,  14'd1310,  -14'd1954,  -14'd313,  -14'd1018,  14'd486,  14'd599,  
-14'd278,  -14'd1662,  -14'd1117,  14'd1208,  14'd1860,  -14'd1089,  -14'd669,  14'd1346,  14'd323,  14'd2512,  14'd1440,  14'd828,  -14'd438,  14'd56,  14'd471,  14'd1763,  

14'd354,  14'd585,  14'd329,  14'd472,  14'd67,  14'd166,  -14'd1518,  14'd72,  14'd197,  -14'd1269,  14'd599,  -14'd174,  -14'd26,  -14'd894,  -14'd87,  14'd550,  
14'd1053,  -14'd85,  -14'd542,  -14'd986,  14'd764,  14'd1405,  14'd74,  -14'd207,  -14'd583,  -14'd485,  -14'd1095,  14'd627,  14'd1345,  -14'd479,  14'd675,  14'd627,  
14'd398,  -14'd329,  14'd114,  14'd671,  14'd190,  14'd875,  -14'd164,  -14'd977,  14'd641,  14'd1062,  -14'd1578,  -14'd1169,  -14'd877,  14'd781,  14'd497,  14'd533,  
-14'd1164,  -14'd275,  -14'd1159,  -14'd361,  -14'd566,  -14'd240,  -14'd393,  -14'd201,  14'd1545,  14'd930,  -14'd229,  -14'd80,  -14'd67,  14'd2018,  14'd1341,  -14'd7,  
-14'd1396,  -14'd689,  -14'd496,  14'd334,  14'd394,  -14'd25,  -14'd1376,  14'd574,  14'd1137,  14'd876,  14'd696,  14'd312,  -14'd1180,  14'd379,  14'd714,  -14'd447,  
14'd374,  14'd109,  -14'd2052,  14'd416,  -14'd646,  -14'd631,  -14'd681,  -14'd1553,  14'd829,  14'd1620,  14'd609,  14'd223,  14'd872,  -14'd1471,  -14'd702,  -14'd257,  
-14'd75,  -14'd9,  -14'd347,  -14'd1066,  14'd840,  14'd280,  -14'd1320,  -14'd349,  -14'd1386,  14'd975,  -14'd391,  -14'd484,  -14'd43,  14'd475,  14'd173,  14'd595,  
-14'd1209,  14'd2271,  14'd572,  -14'd289,  14'd72,  -14'd503,  14'd462,  -14'd862,  14'd1181,  14'd1478,  -14'd403,  14'd1737,  -14'd713,  14'd1376,  -14'd847,  14'd1135,  
14'd129,  -14'd1044,  14'd863,  14'd577,  -14'd260,  14'd130,  -14'd1058,  -14'd292,  -14'd841,  -14'd1627,  -14'd1484,  14'd634,  -14'd34,  14'd1103,  14'd458,  14'd969,  
-14'd582,  14'd859,  14'd1329,  -14'd1341,  -14'd125,  14'd882,  14'd927,  -14'd610,  14'd159,  14'd291,  14'd319,  14'd1128,  -14'd248,  14'd460,  -14'd641,  -14'd614,  
-14'd970,  14'd16,  14'd397,  -14'd468,  -14'd1159,  -14'd9,  14'd141,  -14'd1766,  14'd532,  -14'd618,  14'd706,  14'd17,  -14'd2059,  -14'd1656,  -14'd1363,  14'd830,  
14'd1244,  14'd956,  -14'd667,  14'd211,  -14'd488,  14'd1610,  14'd1003,  -14'd109,  14'd1914,  -14'd163,  -14'd1394,  14'd20,  -14'd438,  14'd426,  -14'd1284,  -14'd722,  
14'd547,  14'd1151,  -14'd1056,  -14'd494,  14'd1115,  -14'd147,  -14'd860,  14'd403,  14'd44,  -14'd435,  -14'd1376,  14'd1690,  14'd1396,  -14'd259,  14'd121,  -14'd1205,  
-14'd509,  14'd54,  14'd745,  14'd671,  -14'd237,  -14'd944,  14'd949,  -14'd1318,  14'd492,  14'd330,  -14'd98,  -14'd125,  14'd4,  14'd461,  -14'd270,  14'd444,  
14'd679,  14'd92,  -14'd1414,  14'd714,  14'd1277,  14'd330,  -14'd463,  -14'd1003,  -14'd782,  14'd118,  -14'd1389,  14'd1095,  14'd748,  -14'd1507,  -14'd772,  -14'd259,  
14'd836,  -14'd1419,  14'd912,  14'd864,  -14'd610,  -14'd106,  14'd1436,  14'd115,  14'd965,  14'd28,  14'd1023,  14'd162,  -14'd662,  14'd602,  14'd44,  14'd132,  
14'd259,  -14'd995,  -14'd247,  14'd764,  14'd315,  14'd1446,  14'd1108,  14'd801,  14'd172,  14'd221,  14'd677,  14'd850,  -14'd460,  14'd573,  14'd839,  14'd64,  
14'd1042,  14'd87,  -14'd918,  14'd1400,  -14'd188,  14'd266,  14'd223,  -14'd123,  -14'd1503,  14'd1067,  14'd104,  14'd40,  14'd742,  -14'd1116,  14'd1038,  -14'd598,  
-14'd317,  -14'd1418,  -14'd1097,  14'd311,  14'd856,  14'd262,  14'd315,  14'd454,  -14'd97,  -14'd484,  14'd1023,  14'd966,  -14'd686,  -14'd1327,  14'd1576,  -14'd587,  
-14'd218,  14'd76,  -14'd1095,  14'd249,  14'd399,  14'd959,  -14'd284,  14'd43,  -14'd685,  14'd1049,  14'd1482,  14'd847,  -14'd395,  -14'd660,  14'd1458,  14'd1525,  
14'd289,  -14'd748,  14'd364,  14'd588,  -14'd645,  -14'd1488,  -14'd913,  14'd451,  -14'd1349,  14'd515,  -14'd115,  -14'd396,  -14'd891,  14'd880,  14'd936,  -14'd1143,  
-14'd768,  -14'd187,  -14'd659,  -14'd1115,  14'd54,  -14'd826,  -14'd957,  14'd112,  -14'd1193,  -14'd256,  14'd1388,  -14'd590,  14'd563,  14'd1807,  14'd394,  14'd809,  
14'd160,  -14'd1646,  -14'd127,  14'd1774,  14'd961,  14'd1313,  -14'd753,  14'd896,  -14'd1934,  -14'd312,  14'd493,  14'd280,  14'd1242,  -14'd619,  14'd811,  14'd820,  
-14'd1046,  14'd25,  -14'd152,  14'd515,  14'd1508,  -14'd149,  14'd561,  14'd663,  14'd754,  14'd1432,  14'd12,  14'd1299,  14'd605,  -14'd360,  -14'd450,  -14'd156,  
14'd326,  14'd2337,  -14'd1217,  14'd1501,  14'd1336,  14'd1396,  14'd217,  -14'd51,  14'd1578,  14'd1802,  14'd552,  14'd252,  14'd196,  -14'd652,  14'd564,  14'd1531,  

14'd273,  14'd582,  -14'd1485,  -14'd304,  14'd225,  -14'd1394,  -14'd1029,  -14'd855,  14'd182,  -14'd69,  14'd259,  14'd891,  -14'd2167,  -14'd1815,  -14'd1127,  14'd4,  
14'd1222,  -14'd977,  -14'd925,  14'd1853,  -14'd303,  14'd190,  -14'd1824,  14'd208,  -14'd434,  14'd458,  14'd974,  -14'd877,  14'd1674,  -14'd686,  14'd17,  14'd1328,  
-14'd630,  14'd515,  -14'd480,  14'd526,  -14'd25,  14'd1475,  -14'd1142,  14'd454,  14'd1528,  14'd1010,  -14'd1363,  14'd795,  14'd1116,  -14'd3394,  -14'd1262,  14'd558,  
-14'd231,  -14'd117,  14'd146,  14'd235,  14'd1014,  14'd204,  -14'd1620,  14'd103,  -14'd1096,  14'd1267,  -14'd99,  14'd1156,  14'd858,  -14'd1458,  -14'd68,  -14'd1258,  
-14'd2067,  -14'd942,  14'd1679,  14'd422,  14'd1116,  14'd60,  -14'd125,  14'd505,  -14'd824,  14'd877,  -14'd350,  -14'd280,  -14'd1113,  -14'd76,  -14'd1246,  -14'd1478,  
14'd58,  -14'd934,  14'd638,  14'd1359,  -14'd699,  14'd1754,  14'd1007,  14'd35,  14'd2310,  14'd878,  14'd351,  14'd624,  14'd761,  14'd24,  -14'd925,  -14'd683,  
-14'd610,  14'd2639,  -14'd675,  14'd52,  -14'd204,  -14'd1049,  -14'd124,  14'd964,  14'd683,  -14'd44,  -14'd555,  14'd645,  14'd726,  -14'd298,  -14'd862,  14'd1229,  
-14'd1678,  14'd636,  14'd188,  -14'd1004,  -14'd284,  14'd1031,  -14'd276,  -14'd882,  -14'd847,  -14'd725,  14'd737,  14'd1083,  14'd756,  -14'd449,  -14'd1168,  14'd2501,  
14'd488,  14'd1040,  14'd209,  -14'd933,  14'd483,  -14'd174,  14'd226,  -14'd491,  14'd1336,  -14'd822,  14'd984,  14'd1391,  -14'd555,  14'd1278,  14'd789,  -14'd154,  
-14'd1278,  -14'd688,  -14'd322,  14'd820,  -14'd160,  -14'd610,  14'd467,  -14'd631,  -14'd710,  -14'd1264,  14'd60,  -14'd844,  -14'd743,  14'd38,  -14'd472,  14'd537,  
14'd1352,  -14'd219,  14'd1493,  14'd342,  14'd2506,  -14'd21,  14'd144,  14'd596,  14'd1060,  14'd377,  -14'd210,  14'd416,  -14'd316,  -14'd487,  14'd586,  14'd836,  
-14'd161,  14'd889,  -14'd593,  -14'd463,  14'd756,  -14'd96,  14'd578,  14'd750,  -14'd2056,  -14'd582,  14'd1376,  14'd469,  14'd83,  -14'd1285,  14'd680,  -14'd1267,  
14'd1944,  -14'd415,  14'd1800,  14'd560,  -14'd758,  -14'd403,  14'd496,  14'd265,  -14'd616,  14'd36,  14'd376,  -14'd696,  -14'd1203,  14'd8,  14'd422,  -14'd1391,  
14'd1488,  14'd613,  14'd711,  -14'd1321,  -14'd477,  -14'd386,  14'd1527,  -14'd1738,  14'd680,  -14'd1414,  -14'd165,  14'd24,  -14'd124,  -14'd47,  -14'd1038,  -14'd805,  
14'd2464,  14'd982,  14'd141,  -14'd611,  -14'd164,  14'd1833,  14'd894,  -14'd230,  14'd581,  -14'd723,  14'd149,  14'd539,  -14'd545,  14'd1796,  -14'd725,  14'd785,  
14'd187,  14'd789,  -14'd54,  14'd725,  14'd729,  -14'd1248,  -14'd702,  14'd373,  -14'd854,  -14'd324,  14'd694,  14'd1487,  14'd585,  14'd608,  14'd1018,  -14'd1220,  
-14'd181,  14'd1809,  -14'd837,  -14'd908,  14'd907,  -14'd138,  -14'd626,  14'd931,  -14'd392,  -14'd3,  -14'd403,  14'd201,  -14'd1127,  -14'd1719,  14'd252,  14'd1269,  
-14'd15,  14'd286,  -14'd1240,  -14'd55,  14'd239,  -14'd838,  -14'd675,  14'd221,  14'd1637,  14'd1180,  -14'd1238,  14'd956,  14'd287,  14'd851,  -14'd563,  14'd444,  
14'd1364,  14'd509,  14'd13,  -14'd562,  -14'd315,  -14'd1506,  14'd120,  -14'd664,  14'd1354,  14'd861,  14'd648,  -14'd917,  -14'd817,  14'd5,  14'd225,  -14'd399,  
-14'd1084,  -14'd1438,  -14'd749,  -14'd235,  -14'd57,  -14'd2304,  14'd989,  -14'd451,  14'd1291,  14'd397,  14'd1005,  -14'd1040,  14'd955,  14'd664,  -14'd1018,  14'd665,  
14'd158,  -14'd148,  -14'd521,  -14'd459,  -14'd1357,  -14'd176,  -14'd1605,  -14'd1351,  -14'd800,  14'd647,  14'd1289,  -14'd389,  14'd336,  14'd1385,  -14'd36,  -14'd104,  
14'd158,  -14'd80,  14'd691,  14'd207,  14'd1304,  14'd188,  14'd379,  14'd53,  14'd534,  14'd529,  -14'd303,  14'd1043,  -14'd413,  -14'd730,  14'd581,  14'd661,  
14'd614,  14'd185,  14'd1085,  -14'd246,  -14'd56,  -14'd38,  14'd480,  14'd1123,  14'd57,  -14'd1151,  -14'd1544,  -14'd1246,  -14'd1323,  -14'd69,  14'd91,  -14'd979,  
-14'd695,  -14'd488,  -14'd1180,  -14'd780,  -14'd428,  14'd856,  -14'd93,  -14'd944,  14'd822,  -14'd670,  -14'd762,  14'd1234,  14'd378,  14'd1029,  14'd1158,  -14'd828,  
-14'd429,  -14'd1087,  14'd509,  14'd583,  -14'd481,  14'd253,  14'd136,  -14'd261,  -14'd1519,  14'd1804,  14'd386,  -14'd1108,  14'd570,  14'd327,  14'd683,  -14'd147,  

-14'd244,  14'd885,  -14'd131,  14'd233,  -14'd1287,  -14'd17,  14'd640,  -14'd98,  -14'd1404,  -14'd218,  14'd2184,  14'd1490,  14'd306,  14'd200,  14'd85,  14'd803,  
-14'd1540,  14'd1271,  -14'd672,  14'd81,  -14'd709,  -14'd6,  14'd480,  14'd59,  -14'd109,  14'd886,  14'd922,  14'd246,  -14'd383,  -14'd1962,  14'd870,  -14'd20,  
-14'd43,  14'd928,  -14'd877,  -14'd1235,  14'd1960,  -14'd399,  14'd333,  14'd835,  14'd559,  14'd677,  14'd896,  -14'd298,  14'd271,  -14'd2889,  -14'd556,  -14'd316,  
-14'd969,  -14'd1766,  14'd301,  14'd983,  -14'd117,  -14'd882,  -14'd665,  14'd1175,  14'd106,  -14'd257,  -14'd166,  14'd1016,  -14'd1284,  14'd313,  -14'd515,  -14'd273,  
-14'd468,  -14'd1280,  14'd1005,  -14'd302,  -14'd1261,  -14'd1047,  -14'd193,  -14'd120,  -14'd78,  14'd269,  -14'd497,  14'd102,  -14'd45,  -14'd534,  -14'd350,  14'd1170,  
14'd431,  14'd1593,  -14'd760,  14'd151,  -14'd376,  14'd400,  -14'd1410,  -14'd393,  -14'd125,  -14'd1517,  14'd754,  -14'd15,  14'd1352,  14'd1070,  14'd855,  14'd1697,  
14'd1251,  14'd184,  -14'd766,  -14'd1159,  14'd532,  -14'd137,  14'd728,  -14'd578,  14'd1189,  -14'd1490,  14'd549,  14'd857,  14'd111,  -14'd203,  14'd1293,  14'd397,  
14'd1123,  14'd848,  -14'd1298,  14'd147,  14'd1148,  -14'd459,  14'd394,  14'd1110,  14'd999,  14'd449,  -14'd713,  14'd2315,  -14'd1214,  -14'd342,  -14'd506,  14'd1140,  
14'd449,  14'd477,  -14'd1587,  -14'd270,  14'd572,  14'd212,  14'd1721,  -14'd470,  -14'd150,  -14'd39,  -14'd1029,  -14'd55,  14'd144,  -14'd386,  14'd233,  14'd354,  
-14'd1539,  -14'd1547,  -14'd838,  14'd452,  14'd359,  -14'd409,  14'd1288,  -14'd39,  14'd457,  -14'd252,  -14'd83,  -14'd307,  14'd148,  14'd870,  -14'd1313,  14'd189,  
-14'd673,  -14'd641,  14'd1217,  14'd558,  -14'd402,  -14'd120,  14'd1215,  -14'd816,  -14'd830,  -14'd353,  -14'd518,  -14'd1000,  -14'd114,  -14'd97,  -14'd665,  -14'd1167,  
14'd1081,  -14'd279,  -14'd1014,  14'd232,  -14'd221,  -14'd1206,  -14'd1183,  -14'd804,  -14'd1164,  -14'd1120,  -14'd52,  -14'd581,  14'd153,  14'd1018,  14'd1438,  14'd98,  
14'd723,  14'd5,  14'd705,  14'd189,  14'd493,  -14'd1001,  -14'd233,  -14'd1187,  -14'd417,  14'd68,  14'd987,  14'd331,  -14'd317,  14'd82,  -14'd567,  -14'd93,  
14'd1041,  -14'd1626,  -14'd443,  -14'd1254,  14'd631,  14'd706,  -14'd1216,  -14'd94,  14'd122,  -14'd43,  14'd587,  -14'd18,  -14'd253,  -14'd164,  14'd443,  14'd285,  
-14'd1558,  -14'd134,  14'd732,  14'd436,  14'd924,  14'd964,  14'd12,  -14'd858,  -14'd10,  14'd1370,  -14'd347,  14'd902,  -14'd692,  14'd30,  -14'd1076,  -14'd47,  
14'd821,  14'd1243,  14'd980,  14'd544,  14'd85,  -14'd46,  -14'd436,  -14'd595,  14'd1298,  14'd872,  -14'd533,  -14'd2342,  14'd354,  -14'd473,  -14'd1090,  -14'd433,  
-14'd1012,  14'd146,  -14'd1385,  -14'd515,  14'd1231,  -14'd614,  14'd522,  14'd87,  -14'd283,  -14'd39,  14'd256,  -14'd377,  14'd421,  -14'd451,  -14'd1556,  -14'd1269,  
14'd190,  -14'd210,  14'd382,  -14'd599,  -14'd1102,  -14'd1051,  14'd193,  14'd1500,  14'd224,  14'd80,  -14'd78,  -14'd1034,  14'd826,  14'd1099,  -14'd543,  14'd999,  
14'd1358,  -14'd356,  14'd832,  14'd956,  14'd129,  14'd163,  -14'd1352,  -14'd976,  -14'd656,  14'd391,  14'd865,  14'd1200,  -14'd976,  14'd1393,  14'd1114,  14'd579,  
14'd1008,  14'd1426,  -14'd1715,  14'd824,  -14'd406,  14'd482,  14'd653,  14'd1326,  -14'd297,  14'd1275,  -14'd194,  -14'd982,  14'd750,  14'd93,  14'd509,  -14'd637,  
14'd742,  14'd343,  -14'd892,  14'd112,  -14'd437,  -14'd983,  14'd496,  -14'd1343,  14'd975,  -14'd312,  14'd841,  14'd3,  14'd82,  -14'd1986,  14'd721,  14'd768,  
14'd1123,  14'd1308,  14'd267,  -14'd1089,  -14'd1771,  -14'd786,  14'd786,  -14'd1842,  14'd2273,  -14'd927,  -14'd1428,  -14'd344,  -14'd662,  -14'd1169,  -14'd1353,  14'd694,  
-14'd1149,  14'd458,  14'd1041,  -14'd843,  -14'd518,  14'd476,  14'd28,  -14'd305,  14'd2089,  14'd2811,  -14'd1483,  14'd599,  14'd30,  14'd2606,  14'd876,  -14'd162,  
14'd1027,  -14'd1007,  14'd375,  -14'd107,  -14'd340,  14'd41,  14'd784,  14'd1121,  14'd1418,  -14'd800,  -14'd970,  14'd1398,  -14'd48,  14'd1585,  -14'd1166,  -14'd658,  
-14'd785,  14'd1321,  14'd1798,  14'd1419,  14'd383,  -14'd407,  14'd1656,  14'd1406,  14'd1399,  -14'd361,  -14'd1359,  -14'd110,  14'd827,  14'd340,  14'd374,  14'd132,  

-14'd824,  -14'd578,  -14'd839,  14'd650,  14'd972,  -14'd619,  -14'd2893,  14'd446,  -14'd762,  -14'd262,  -14'd1078,  -14'd125,  14'd663,  -14'd388,  14'd1441,  14'd1086,  
-14'd718,  -14'd362,  -14'd330,  14'd341,  -14'd586,  -14'd950,  -14'd91,  14'd1595,  -14'd332,  14'd1479,  -14'd459,  -14'd312,  14'd311,  -14'd1699,  -14'd513,  -14'd92,  
-14'd848,  14'd969,  14'd555,  14'd1938,  14'd110,  -14'd940,  -14'd1269,  14'd1526,  -14'd1007,  -14'd663,  -14'd1443,  14'd420,  14'd398,  -14'd2467,  -14'd167,  14'd1453,  
14'd500,  -14'd609,  -14'd639,  14'd946,  -14'd464,  14'd993,  -14'd550,  14'd539,  -14'd61,  14'd840,  14'd1001,  14'd333,  14'd1161,  -14'd1200,  -14'd176,  14'd2285,  
-14'd337,  -14'd1741,  14'd332,  14'd97,  14'd49,  14'd169,  14'd1203,  -14'd873,  14'd837,  14'd2140,  14'd334,  14'd682,  14'd698,  -14'd489,  -14'd396,  14'd199,  
-14'd1042,  14'd607,  14'd96,  14'd1004,  14'd1117,  14'd117,  -14'd1399,  -14'd1001,  14'd650,  14'd467,  -14'd819,  14'd1537,  14'd1347,  -14'd1497,  -14'd1840,  14'd965,  
-14'd588,  -14'd136,  -14'd497,  -14'd354,  14'd526,  14'd85,  14'd630,  -14'd83,  -14'd53,  -14'd940,  14'd386,  -14'd796,  14'd870,  -14'd1453,  -14'd1352,  14'd413,  
-14'd25,  14'd253,  -14'd797,  14'd680,  14'd285,  -14'd149,  14'd563,  -14'd360,  -14'd1653,  14'd1458,  14'd709,  -14'd759,  14'd711,  14'd2087,  14'd100,  14'd822,  
14'd207,  14'd337,  14'd2108,  -14'd850,  -14'd121,  14'd1047,  14'd415,  -14'd361,  -14'd744,  14'd284,  14'd288,  14'd1082,  14'd116,  14'd697,  14'd962,  14'd2310,  
14'd4,  -14'd156,  -14'd1022,  14'd770,  14'd25,  14'd676,  14'd1373,  14'd780,  14'd109,  -14'd406,  -14'd414,  14'd47,  -14'd57,  14'd833,  14'd265,  -14'd465,  
-14'd1091,  14'd1086,  -14'd1310,  14'd430,  -14'd296,  -14'd221,  14'd124,  14'd843,  14'd1712,  -14'd1569,  14'd280,  14'd130,  -14'd603,  -14'd1448,  -14'd986,  14'd555,  
14'd313,  -14'd1460,  -14'd669,  -14'd2065,  14'd1536,  14'd0,  14'd262,  -14'd283,  14'd190,  -14'd456,  -14'd26,  -14'd630,  14'd1209,  -14'd260,  14'd522,  14'd277,  
-14'd552,  -14'd731,  14'd1381,  14'd649,  14'd772,  14'd39,  -14'd636,  -14'd1535,  -14'd728,  -14'd256,  -14'd1206,  14'd44,  -14'd838,  14'd785,  14'd786,  -14'd619,  
14'd812,  14'd1273,  14'd488,  -14'd631,  14'd1628,  14'd1374,  14'd735,  14'd1457,  14'd932,  14'd1166,  14'd222,  14'd716,  14'd1295,  14'd420,  -14'd276,  14'd21,  
14'd1692,  -14'd408,  14'd1496,  -14'd5,  14'd823,  14'd1107,  14'd1043,  14'd307,  -14'd1252,  -14'd1183,  -14'd253,  14'd1084,  14'd939,  14'd61,  14'd897,  14'd555,  
14'd359,  14'd148,  -14'd161,  14'd862,  -14'd899,  -14'd478,  14'd429,  14'd719,  14'd586,  14'd352,  -14'd785,  14'd554,  -14'd1206,  -14'd483,  14'd459,  14'd218,  
14'd1431,  14'd41,  -14'd38,  -14'd592,  -14'd371,  14'd638,  -14'd979,  14'd15,  14'd785,  14'd413,  14'd274,  -14'd401,  14'd19,  14'd613,  -14'd4,  -14'd743,  
-14'd692,  14'd246,  14'd607,  14'd1114,  14'd79,  -14'd1084,  14'd147,  14'd1158,  14'd143,  -14'd1392,  14'd1148,  -14'd387,  -14'd226,  -14'd339,  -14'd33,  -14'd436,  
-14'd1474,  -14'd1256,  14'd124,  14'd99,  -14'd576,  -14'd678,  14'd1045,  -14'd516,  -14'd1008,  -14'd1111,  14'd1578,  14'd967,  14'd835,  14'd43,  14'd1269,  -14'd274,  
14'd636,  -14'd162,  -14'd280,  -14'd1574,  14'd531,  14'd252,  14'd806,  -14'd649,  -14'd1358,  -14'd391,  14'd1160,  -14'd98,  -14'd141,  -14'd1066,  -14'd479,  14'd651,  
-14'd345,  14'd154,  -14'd33,  -14'd358,  14'd15,  -14'd740,  -14'd475,  -14'd71,  -14'd1256,  14'd28,  -14'd126,  -14'd149,  -14'd894,  -14'd936,  14'd1340,  14'd430,  
-14'd351,  14'd493,  -14'd526,  -14'd245,  -14'd273,  -14'd1441,  -14'd36,  -14'd1573,  14'd600,  -14'd1368,  -14'd218,  14'd391,  14'd770,  14'd383,  -14'd1125,  14'd972,  
14'd126,  14'd497,  14'd474,  -14'd1515,  -14'd1358,  -14'd1579,  -14'd185,  14'd803,  -14'd84,  14'd1679,  -14'd1631,  14'd746,  -14'd1080,  14'd423,  -14'd1324,  -14'd53,  
-14'd662,  14'd621,  14'd809,  -14'd658,  14'd646,  -14'd202,  14'd861,  -14'd509,  -14'd1251,  -14'd228,  14'd70,  14'd400,  -14'd1165,  -14'd1211,  14'd484,  -14'd1028,  
14'd413,  14'd825,  14'd12,  -14'd1593,  14'd31,  -14'd1772,  -14'd567,  -14'd224,  -14'd1201,  -14'd685,  14'd546,  -14'd2268,  -14'd915,  -14'd624,  -14'd1754,  -14'd358,  

-14'd828,  14'd1165,  -14'd219,  14'd308,  14'd826,  14'd854,  -14'd788,  -14'd90,  14'd1508,  14'd330,  14'd260,  -14'd1155,  -14'd289,  14'd625,  -14'd499,  -14'd766,  
-14'd1059,  -14'd423,  14'd1787,  14'd1326,  14'd577,  14'd470,  14'd586,  14'd86,  -14'd393,  -14'd403,  -14'd666,  14'd17,  14'd1576,  14'd395,  14'd1518,  14'd1516,  
14'd759,  -14'd1270,  14'd918,  -14'd821,  -14'd112,  14'd482,  14'd1515,  14'd431,  14'd495,  14'd1285,  14'd949,  14'd899,  -14'd367,  14'd1412,  14'd1098,  -14'd781,  
14'd797,  -14'd452,  -14'd302,  14'd1235,  -14'd724,  -14'd207,  14'd542,  -14'd1120,  14'd1776,  14'd181,  14'd515,  -14'd906,  -14'd335,  14'd1579,  -14'd2080,  -14'd559,  
14'd430,  -14'd330,  -14'd1147,  -14'd1536,  14'd1058,  -14'd1149,  14'd1492,  14'd269,  14'd61,  -14'd669,  14'd993,  -14'd409,  14'd579,  -14'd709,  -14'd1000,  -14'd569,  
-14'd1457,  -14'd791,  -14'd468,  -14'd1709,  14'd1366,  -14'd1077,  14'd407,  14'd833,  -14'd856,  14'd361,  14'd300,  -14'd1706,  -14'd935,  -14'd1216,  14'd150,  14'd116,  
-14'd752,  -14'd718,  14'd158,  14'd508,  -14'd305,  -14'd881,  -14'd2730,  -14'd512,  -14'd1271,  14'd1208,  -14'd612,  -14'd1303,  -14'd695,  -14'd2190,  14'd47,  14'd33,  
14'd909,  -14'd2590,  14'd1593,  14'd498,  -14'd87,  14'd1423,  14'd131,  14'd33,  -14'd3111,  14'd86,  14'd181,  -14'd367,  -14'd629,  14'd365,  14'd786,  14'd355,  
14'd1729,  -14'd803,  14'd1396,  14'd814,  14'd170,  -14'd667,  14'd1093,  14'd2137,  -14'd1745,  -14'd290,  14'd957,  -14'd1159,  -14'd607,  14'd1154,  14'd138,  -14'd119,  
14'd2440,  -14'd1048,  14'd867,  14'd1077,  -14'd607,  -14'd125,  -14'd685,  -14'd320,  14'd813,  14'd917,  14'd581,  -14'd1265,  -14'd270,  14'd402,  -14'd1356,  -14'd28,  
-14'd1454,  -14'd519,  -14'd2027,  -14'd8,  14'd804,  -14'd1175,  -14'd481,  14'd485,  14'd1000,  14'd161,  -14'd299,  -14'd2468,  14'd292,  -14'd2597,  -14'd663,  -14'd1180,  
-14'd94,  -14'd705,  -14'd557,  14'd488,  -14'd1620,  14'd138,  -14'd1620,  -14'd511,  14'd298,  14'd343,  14'd205,  14'd302,  -14'd1619,  -14'd144,  14'd762,  14'd663,  
14'd1834,  14'd782,  14'd1270,  14'd225,  -14'd1738,  14'd35,  -14'd1569,  14'd513,  -14'd514,  14'd1667,  14'd1002,  -14'd460,  14'd522,  -14'd212,  14'd2035,  14'd762,  
14'd699,  -14'd889,  14'd312,  14'd267,  -14'd228,  14'd175,  -14'd680,  14'd890,  -14'd1084,  14'd1090,  -14'd565,  -14'd1296,  14'd1996,  -14'd1034,  -14'd836,  14'd488,  
-14'd1026,  -14'd760,  -14'd99,  14'd770,  -14'd1183,  -14'd1127,  14'd646,  14'd516,  14'd1087,  -14'd260,  14'd872,  -14'd197,  -14'd249,  14'd163,  -14'd631,  -14'd34,  
-14'd2038,  -14'd91,  -14'd1015,  14'd358,  14'd199,  14'd410,  14'd108,  14'd575,  14'd532,  14'd923,  14'd627,  -14'd1784,  -14'd1324,  14'd778,  14'd267,  -14'd655,  
14'd742,  14'd999,  -14'd507,  -14'd217,  -14'd937,  14'd1227,  14'd395,  -14'd98,  -14'd1057,  14'd461,  14'd291,  -14'd177,  14'd453,  -14'd223,  14'd434,  -14'd592,  
14'd612,  -14'd28,  -14'd1188,  14'd711,  -14'd557,  -14'd71,  14'd499,  14'd732,  -14'd169,  14'd351,  14'd644,  14'd225,  14'd1225,  -14'd1504,  14'd432,  14'd676,  
-14'd15,  -14'd597,  14'd1519,  14'd407,  -14'd983,  -14'd617,  -14'd917,  -14'd372,  -14'd733,  14'd231,  14'd924,  14'd128,  -14'd755,  -14'd212,  14'd28,  14'd41,  
-14'd816,  -14'd270,  14'd11,  -14'd236,  14'd300,  -14'd417,  14'd241,  14'd1089,  -14'd745,  14'd1275,  -14'd126,  -14'd401,  -14'd96,  14'd683,  -14'd766,  -14'd251,  
14'd425,  14'd1476,  -14'd444,  14'd881,  -14'd205,  14'd767,  14'd1038,  -14'd450,  14'd934,  -14'd258,  -14'd702,  14'd1265,  14'd332,  -14'd549,  14'd436,  -14'd170,  
14'd56,  14'd1060,  14'd340,  -14'd126,  14'd340,  -14'd85,  14'd507,  14'd410,  -14'd595,  -14'd274,  -14'd1095,  14'd108,  14'd346,  14'd949,  14'd1004,  -14'd652,  
14'd715,  -14'd417,  14'd489,  -14'd677,  14'd715,  14'd591,  14'd527,  -14'd555,  14'd703,  14'd1100,  14'd763,  -14'd162,  -14'd649,  -14'd890,  14'd834,  14'd721,  
-14'd468,  14'd540,  -14'd83,  -14'd752,  -14'd952,  -14'd1615,  14'd1053,  -14'd1022,  -14'd951,  -14'd674,  14'd284,  14'd241,  -14'd902,  14'd1763,  14'd528,  14'd553,  
14'd639,  14'd1412,  -14'd80,  14'd709,  14'd515,  -14'd1339,  -14'd877,  -14'd588,  14'd1477,  -14'd832,  14'd529,  -14'd255,  -14'd1827,  14'd1282,  -14'd904,  -14'd92,  

-14'd1339,  14'd830,  -14'd570,  -14'd813,  -14'd393,  14'd3,  -14'd346,  -14'd1319,  -14'd926,  -14'd1404,  -14'd2130,  -14'd998,  -14'd681,  -14'd1296,  -14'd870,  -14'd879,  
-14'd1123,  14'd933,  -14'd252,  14'd1097,  -14'd269,  14'd1641,  14'd381,  14'd344,  14'd714,  -14'd260,  -14'd2367,  14'd275,  -14'd1052,  14'd505,  14'd116,  14'd405,  
14'd935,  -14'd132,  -14'd509,  14'd175,  14'd1824,  14'd1291,  14'd995,  -14'd1152,  -14'd1558,  -14'd956,  14'd931,  14'd693,  -14'd1119,  -14'd731,  14'd749,  -14'd1480,  
-14'd911,  -14'd391,  -14'd76,  14'd1207,  -14'd96,  14'd1236,  -14'd767,  -14'd230,  -14'd343,  -14'd456,  14'd685,  -14'd628,  14'd1538,  14'd2527,  -14'd656,  -14'd1337,  
-14'd917,  -14'd1471,  -14'd437,  14'd1157,  14'd1444,  -14'd316,  14'd451,  14'd82,  -14'd1405,  14'd726,  -14'd610,  -14'd1373,  -14'd779,  -14'd396,  14'd606,  -14'd1575,  
-14'd925,  -14'd553,  -14'd1663,  14'd302,  14'd1724,  -14'd1708,  -14'd355,  -14'd1618,  14'd322,  -14'd488,  -14'd133,  14'd686,  -14'd377,  -14'd121,  -14'd1492,  -14'd1754,  
14'd815,  -14'd217,  14'd702,  -14'd1618,  14'd1101,  -14'd611,  -14'd417,  -14'd712,  -14'd965,  14'd442,  -14'd1145,  -14'd1789,  -14'd1926,  -14'd1011,  -14'd415,  -14'd1590,  
14'd693,  14'd1256,  14'd848,  14'd40,  -14'd1875,  14'd145,  -14'd179,  14'd494,  14'd924,  14'd674,  -14'd377,  -14'd774,  -14'd588,  14'd631,  14'd930,  -14'd1241,  
14'd55,  14'd26,  14'd1117,  14'd295,  -14'd205,  -14'd716,  14'd1274,  -14'd576,  -14'd631,  -14'd589,  14'd893,  14'd1211,  14'd394,  14'd2468,  14'd753,  14'd738,  
-14'd698,  14'd509,  14'd602,  -14'd553,  -14'd35,  -14'd373,  14'd622,  -14'd1159,  14'd368,  -14'd341,  -14'd89,  14'd240,  -14'd573,  -14'd246,  -14'd1305,  -14'd1029,  
-14'd1374,  -14'd1186,  -14'd35,  14'd642,  14'd153,  -14'd642,  -14'd138,  14'd231,  14'd1405,  -14'd589,  14'd499,  -14'd441,  -14'd286,  14'd625,  -14'd142,  -14'd1324,  
-14'd338,  -14'd1108,  14'd99,  14'd902,  14'd688,  14'd1524,  14'd323,  -14'd267,  14'd894,  -14'd267,  -14'd297,  -14'd809,  14'd236,  -14'd630,  14'd365,  14'd461,  
14'd916,  14'd111,  14'd804,  -14'd789,  14'd654,  14'd1617,  -14'd80,  14'd1125,  14'd1188,  -14'd235,  -14'd1173,  14'd897,  -14'd1,  14'd250,  14'd830,  -14'd1283,  
14'd577,  -14'd500,  14'd485,  -14'd177,  -14'd25,  14'd529,  14'd655,  14'd563,  14'd1158,  14'd210,  -14'd730,  -14'd95,  14'd962,  14'd1040,  14'd579,  -14'd783,  
14'd839,  14'd1274,  -14'd134,  14'd476,  14'd222,  -14'd1906,  -14'd777,  -14'd33,  -14'd1427,  -14'd1990,  14'd268,  -14'd915,  -14'd531,  -14'd808,  -14'd34,  14'd125,  
14'd795,  -14'd380,  14'd832,  14'd258,  -14'd592,  -14'd982,  14'd1140,  -14'd1122,  14'd314,  -14'd1969,  14'd2269,  14'd1256,  14'd474,  -14'd507,  -14'd337,  14'd649,  
14'd449,  -14'd385,  -14'd14,  -14'd946,  -14'd2435,  14'd226,  14'd1112,  -14'd105,  14'd409,  14'd355,  14'd1070,  -14'd1191,  14'd839,  14'd1238,  14'd395,  14'd1592,  
14'd786,  -14'd810,  -14'd862,  14'd959,  -14'd846,  14'd1168,  14'd276,  14'd1817,  14'd1108,  -14'd783,  14'd1138,  -14'd910,  14'd484,  14'd1200,  14'd1297,  14'd386,  
-14'd343,  -14'd752,  -14'd937,  -14'd50,  -14'd365,  14'd232,  14'd708,  14'd1390,  -14'd743,  14'd947,  -14'd75,  14'd137,  -14'd312,  14'd1377,  -14'd337,  -14'd254,  
14'd1113,  14'd639,  -14'd384,  14'd325,  -14'd2461,  -14'd728,  -14'd2079,  -14'd1260,  -14'd2127,  -14'd2313,  14'd432,  14'd654,  -14'd1657,  14'd1718,  -14'd415,  -14'd774,  
14'd269,  -14'd1868,  14'd172,  -14'd1093,  -14'd1212,  14'd268,  14'd1558,  -14'd553,  14'd276,  14'd389,  14'd508,  -14'd6,  -14'd890,  14'd947,  14'd20,  -14'd759,  
14'd901,  14'd390,  -14'd88,  -14'd1349,  14'd343,  14'd470,  14'd1722,  -14'd1424,  14'd1978,  14'd1500,  14'd46,  -14'd159,  -14'd1314,  14'd17,  -14'd510,  14'd346,  
14'd124,  -14'd529,  14'd2159,  -14'd1282,  14'd875,  -14'd608,  -14'd260,  14'd650,  14'd1018,  14'd997,  -14'd1220,  14'd204,  -14'd1019,  14'd1104,  14'd860,  -14'd1002,  
-14'd2304,  -14'd1182,  -14'd420,  14'd787,  14'd1447,  -14'd381,  14'd1225,  -14'd153,  14'd89,  14'd424,  -14'd681,  -14'd1231,  14'd99,  -14'd331,  14'd148,  -14'd1030,  
14'd11,  14'd517,  14'd1662,  14'd427,  -14'd24,  14'd369,  -14'd824,  14'd249,  14'd75,  14'd709,  -14'd1253,  14'd543,  14'd1574,  14'd164,  -14'd796,  14'd222,  

-14'd916,  -14'd426,  -14'd1187,  14'd1260,  14'd1078,  -14'd728,  14'd352,  14'd815,  -14'd1333,  -14'd978,  14'd1481,  -14'd1947,  14'd530,  -14'd1239,  -14'd853,  14'd41,  
14'd225,  -14'd539,  -14'd834,  14'd1200,  14'd331,  14'd835,  -14'd379,  14'd553,  14'd185,  -14'd548,  -14'd1286,  -14'd68,  14'd1345,  -14'd2103,  -14'd557,  -14'd875,  
-14'd782,  -14'd1065,  -14'd1259,  14'd558,  -14'd15,  -14'd489,  -14'd1582,  -14'd98,  -14'd942,  -14'd598,  14'd683,  -14'd1605,  -14'd507,  -14'd1298,  -14'd871,  14'd464,  
-14'd862,  -14'd2130,  14'd1005,  14'd1033,  14'd784,  -14'd23,  14'd259,  -14'd594,  -14'd575,  14'd1286,  14'd402,  -14'd191,  -14'd480,  -14'd803,  14'd1328,  14'd965,  
-14'd905,  -14'd1751,  14'd621,  -14'd224,  -14'd247,  -14'd181,  -14'd115,  -14'd1021,  14'd1108,  -14'd978,  -14'd213,  -14'd21,  -14'd1543,  14'd56,  -14'd37,  -14'd236,  
-14'd862,  14'd192,  -14'd1817,  14'd30,  -14'd1251,  -14'd1616,  14'd43,  -14'd659,  -14'd207,  -14'd470,  14'd1949,  -14'd647,  14'd434,  14'd126,  -14'd826,  -14'd1450,  
-14'd395,  -14'd1242,  -14'd569,  14'd385,  14'd775,  -14'd1536,  14'd645,  -14'd1249,  -14'd352,  14'd574,  -14'd378,  14'd1745,  -14'd812,  -14'd1710,  14'd904,  14'd363,  
-14'd175,  14'd551,  -14'd390,  14'd164,  14'd1445,  14'd599,  14'd477,  -14'd209,  14'd346,  14'd877,  14'd433,  14'd1398,  14'd869,  14'd45,  14'd389,  14'd937,  
14'd1018,  -14'd879,  -14'd1379,  -14'd343,  14'd1724,  14'd276,  -14'd53,  14'd925,  -14'd253,  14'd959,  14'd6,  14'd1811,  14'd113,  14'd185,  -14'd117,  14'd199,  
-14'd1145,  14'd1070,  14'd1166,  14'd1623,  -14'd78,  14'd166,  14'd1686,  14'd303,  14'd520,  14'd1538,  14'd298,  14'd1209,  -14'd292,  -14'd452,  14'd1254,  14'd203,  
-14'd860,  14'd920,  14'd1170,  14'd805,  -14'd831,  14'd166,  -14'd829,  -14'd658,  14'd248,  -14'd674,  14'd219,  -14'd484,  -14'd949,  -14'd1482,  -14'd1288,  -14'd995,  
14'd27,  -14'd125,  -14'd177,  -14'd603,  -14'd676,  -14'd185,  -14'd1426,  14'd246,  -14'd115,  14'd413,  -14'd1357,  14'd382,  -14'd1017,  -14'd2227,  -14'd486,  -14'd179,  
14'd1599,  -14'd1548,  -14'd525,  -14'd844,  -14'd495,  -14'd1900,  -14'd786,  -14'd27,  14'd356,  14'd763,  14'd358,  -14'd257,  -14'd309,  -14'd842,  14'd1256,  14'd955,  
-14'd624,  -14'd241,  14'd492,  -14'd882,  14'd887,  14'd500,  14'd183,  14'd1037,  -14'd955,  14'd179,  14'd994,  -14'd269,  14'd479,  -14'd884,  -14'd73,  14'd615,  
-14'd156,  -14'd723,  -14'd38,  14'd1080,  14'd1134,  14'd91,  -14'd437,  14'd1168,  14'd95,  14'd31,  -14'd336,  14'd1060,  -14'd894,  14'd162,  14'd1,  -14'd69,  
-14'd844,  -14'd636,  14'd190,  -14'd82,  -14'd1045,  14'd1040,  -14'd2044,  14'd760,  14'd1178,  14'd53,  -14'd683,  -14'd1096,  14'd1393,  14'd1036,  -14'd1051,  14'd379,  
-14'd238,  -14'd1913,  -14'd1438,  14'd531,  -14'd47,  -14'd642,  -14'd1091,  14'd1335,  -14'd1332,  14'd863,  14'd1071,  14'd586,  14'd682,  -14'd226,  -14'd64,  14'd662,  
-14'd1439,  14'd539,  -14'd553,  -14'd653,  14'd1023,  -14'd1298,  -14'd127,  14'd738,  -14'd749,  -14'd948,  14'd138,  -14'd761,  14'd775,  -14'd852,  14'd1022,  -14'd900,  
14'd595,  14'd820,  14'd681,  14'd96,  14'd1336,  14'd531,  -14'd497,  -14'd455,  -14'd420,  14'd852,  -14'd434,  14'd382,  -14'd592,  14'd204,  14'd538,  14'd610,  
14'd223,  -14'd270,  14'd954,  -14'd624,  -14'd94,  -14'd321,  14'd916,  14'd43,  -14'd708,  14'd1155,  14'd951,  -14'd814,  14'd1557,  -14'd430,  14'd564,  -14'd166,  
-14'd763,  -14'd71,  14'd458,  -14'd237,  14'd40,  14'd447,  -14'd1139,  14'd307,  14'd285,  14'd448,  -14'd96,  -14'd406,  14'd577,  14'd225,  14'd1166,  -14'd449,  
14'd10,  14'd118,  14'd111,  14'd795,  14'd906,  -14'd120,  14'd1211,  -14'd1045,  -14'd1789,  -14'd1075,  -14'd22,  14'd1352,  14'd315,  -14'd1156,  -14'd734,  14'd3,  
-14'd131,  14'd141,  14'd200,  14'd167,  14'd1204,  14'd357,  -14'd72,  -14'd1104,  -14'd182,  14'd654,  -14'd494,  14'd1604,  14'd1423,  -14'd893,  -14'd92,  14'd1189,  
14'd959,  14'd1540,  -14'd761,  -14'd695,  14'd572,  14'd396,  14'd252,  -14'd1305,  14'd1000,  -14'd46,  -14'd190,  -14'd788,  14'd789,  -14'd408,  -14'd725,  14'd1275,  
14'd1550,  14'd2367,  14'd843,  -14'd169,  14'd1146,  14'd1005,  -14'd260,  14'd1315,  14'd2127,  14'd3005,  -14'd618,  14'd1485,  -14'd1324,  14'd1588,  14'd430,  14'd807,  

14'd337,  14'd288,  14'd1768,  14'd337,  -14'd255,  14'd301,  14'd825,  -14'd400,  14'd633,  14'd942,  -14'd388,  -14'd359,  14'd322,  14'd536,  -14'd1244,  14'd710,  
-14'd122,  -14'd321,  14'd407,  -14'd617,  -14'd784,  14'd29,  14'd504,  -14'd486,  -14'd750,  -14'd209,  14'd1445,  14'd35,  -14'd674,  14'd2494,  -14'd1544,  14'd215,  
-14'd515,  -14'd1869,  14'd1124,  -14'd414,  -14'd1743,  -14'd428,  14'd939,  14'd807,  -14'd377,  14'd898,  14'd1224,  -14'd896,  14'd1407,  14'd1617,  -14'd866,  -14'd1416,  
14'd1374,  14'd1688,  -14'd563,  14'd135,  14'd399,  -14'd544,  14'd733,  14'd716,  -14'd10,  -14'd272,  14'd1116,  14'd1478,  14'd90,  -14'd170,  -14'd756,  -14'd410,  
14'd2801,  14'd2057,  -14'd877,  14'd803,  -14'd512,  14'd1571,  -14'd197,  14'd365,  -14'd1068,  14'd266,  -14'd58,  14'd1387,  14'd918,  14'd310,  14'd603,  14'd154,  
14'd206,  14'd84,  14'd126,  14'd588,  -14'd605,  14'd1326,  14'd1463,  14'd34,  14'd299,  -14'd289,  14'd130,  14'd23,  -14'd222,  14'd985,  14'd1420,  -14'd422,  
14'd404,  -14'd1525,  -14'd417,  14'd681,  -14'd5,  14'd662,  14'd767,  14'd549,  14'd298,  -14'd884,  14'd2123,  14'd67,  -14'd613,  14'd84,  14'd866,  -14'd1389,  
-14'd1168,  -14'd453,  -14'd461,  -14'd348,  -14'd2161,  -14'd34,  -14'd338,  -14'd1361,  14'd505,  14'd72,  14'd748,  -14'd2046,  14'd879,  14'd503,  -14'd509,  -14'd1068,  
-14'd222,  -14'd264,  -14'd1767,  14'd812,  14'd619,  -14'd1373,  -14'd719,  14'd462,  -14'd30,  14'd302,  14'd561,  14'd193,  14'd580,  -14'd26,  -14'd688,  -14'd654,  
14'd360,  -14'd1896,  -14'd1244,  14'd502,  14'd88,  14'd1152,  -14'd1615,  -14'd847,  14'd603,  14'd294,  -14'd371,  14'd804,  -14'd88,  -14'd238,  -14'd1055,  14'd1872,  
-14'd826,  14'd608,  14'd497,  14'd915,  -14'd11,  14'd691,  14'd474,  14'd593,  -14'd1013,  -14'd942,  -14'd63,  14'd290,  14'd1513,  14'd836,  14'd1535,  14'd358,  
14'd561,  -14'd1031,  14'd261,  14'd200,  14'd1347,  14'd209,  -14'd125,  14'd1188,  14'd333,  -14'd671,  14'd2077,  14'd493,  -14'd137,  -14'd1208,  -14'd184,  14'd648,  
-14'd574,  -14'd481,  -14'd914,  14'd883,  -14'd513,  -14'd1350,  14'd8,  -14'd415,  -14'd517,  14'd1386,  14'd644,  -14'd306,  -14'd804,  14'd64,  -14'd1886,  -14'd209,  
-14'd746,  14'd181,  -14'd908,  14'd1092,  14'd1733,  14'd285,  14'd280,  -14'd651,  14'd158,  14'd902,  14'd460,  14'd78,  -14'd569,  14'd815,  14'd821,  14'd14,  
-14'd1490,  -14'd302,  14'd677,  14'd1200,  -14'd141,  -14'd1256,  -14'd1353,  -14'd636,  14'd512,  14'd1647,  14'd178,  -14'd1032,  -14'd954,  -14'd317,  14'd442,  14'd322,  
-14'd419,  14'd766,  -14'd832,  14'd1099,  14'd1025,  -14'd600,  14'd291,  14'd1289,  14'd106,  -14'd62,  -14'd14,  -14'd1732,  14'd1261,  -14'd212,  -14'd234,  14'd1859,  
-14'd1859,  14'd1633,  -14'd323,  14'd709,  14'd639,  -14'd212,  14'd58,  -14'd7,  -14'd384,  -14'd1123,  -14'd1727,  14'd1075,  14'd711,  -14'd1494,  -14'd821,  14'd287,  
-14'd1174,  -14'd581,  -14'd1180,  -14'd733,  14'd1015,  14'd762,  -14'd289,  -14'd296,  14'd230,  14'd802,  14'd440,  14'd1444,  14'd778,  14'd1621,  -14'd42,  14'd1453,  
14'd182,  -14'd1526,  14'd122,  -14'd550,  14'd1164,  14'd4,  14'd350,  14'd183,  14'd645,  14'd174,  14'd901,  14'd1450,  14'd307,  14'd124,  -14'd360,  14'd1443,  
-14'd923,  14'd5,  14'd1565,  -14'd552,  14'd1136,  14'd91,  14'd1444,  -14'd100,  14'd118,  14'd675,  14'd185,  -14'd592,  -14'd637,  14'd308,  -14'd783,  14'd257,  
14'd799,  -14'd423,  -14'd1331,  -14'd1442,  14'd606,  -14'd387,  14'd1227,  -14'd698,  14'd726,  14'd311,  14'd306,  14'd976,  -14'd684,  -14'd1932,  -14'd649,  14'd334,  
14'd449,  14'd1242,  -14'd377,  -14'd1239,  14'd1567,  14'd462,  14'd1584,  14'd637,  14'd331,  -14'd878,  -14'd912,  -14'd270,  14'd357,  -14'd552,  -14'd361,  14'd225,  
-14'd612,  14'd151,  14'd675,  -14'd344,  14'd1111,  -14'd1751,  14'd950,  -14'd467,  14'd821,  14'd828,  -14'd468,  14'd588,  14'd233,  14'd119,  14'd1189,  14'd148,  
14'd1133,  -14'd334,  14'd1524,  -14'd99,  14'd74,  -14'd1314,  -14'd617,  14'd184,  -14'd104,  14'd1032,  14'd764,  -14'd743,  14'd761,  14'd1878,  -14'd419,  -14'd190,  
14'd1159,  -14'd178,  -14'd676,  -14'd322,  -14'd383,  14'd1860,  14'd193,  14'd780,  -14'd199,  -14'd45,  -14'd680,  14'd506,  -14'd644,  14'd877,  14'd1887,  -14'd522,  

-14'd1654,  -14'd1840,  -14'd648,  -14'd628,  14'd499,  -14'd453,  -14'd1531,  -14'd379,  14'd315,  14'd377,  -14'd1402,  -14'd802,  -14'd2042,  -14'd1518,  14'd516,  -14'd227,  
14'd718,  -14'd353,  14'd650,  -14'd521,  -14'd245,  14'd1155,  14'd121,  -14'd209,  -14'd821,  -14'd198,  -14'd1312,  14'd1485,  14'd825,  14'd1081,  -14'd1000,  -14'd77,  
14'd903,  -14'd665,  14'd616,  14'd669,  14'd472,  -14'd332,  -14'd292,  -14'd709,  14'd119,  -14'd1375,  -14'd695,  14'd1284,  -14'd17,  -14'd133,  -14'd103,  -14'd1165,  
14'd1381,  -14'd1632,  -14'd836,  14'd112,  -14'd295,  14'd203,  14'd1520,  -14'd340,  -14'd148,  14'd1505,  14'd107,  14'd151,  14'd50,  14'd2885,  14'd233,  -14'd1430,  
-14'd1834,  14'd1020,  14'd1027,  -14'd152,  14'd351,  -14'd672,  -14'd923,  14'd34,  14'd93,  14'd1034,  14'd269,  -14'd796,  -14'd1576,  -14'd258,  14'd329,  -14'd1228,  
14'd802,  14'd1167,  -14'd298,  -14'd277,  14'd637,  14'd1167,  14'd691,  -14'd1792,  14'd1413,  -14'd465,  14'd669,  14'd1060,  -14'd1783,  14'd630,  -14'd552,  14'd124,  
-14'd588,  14'd1312,  14'd742,  -14'd554,  -14'd894,  14'd1536,  -14'd1085,  14'd863,  -14'd748,  14'd1416,  -14'd1221,  14'd266,  14'd969,  14'd644,  -14'd244,  -14'd748,  
14'd1341,  -14'd1374,  14'd700,  14'd38,  -14'd839,  14'd1570,  14'd1143,  14'd956,  -14'd1776,  14'd110,  -14'd367,  14'd1073,  -14'd976,  -14'd179,  -14'd55,  -14'd494,  
14'd1054,  14'd805,  14'd1973,  14'd535,  14'd1299,  14'd36,  14'd1146,  14'd125,  -14'd754,  -14'd1037,  14'd45,  14'd346,  14'd272,  14'd1043,  -14'd445,  -14'd527,  
14'd723,  14'd405,  14'd1605,  14'd648,  -14'd385,  -14'd679,  14'd91,  14'd846,  -14'd770,  -14'd1653,  14'd669,  14'd656,  14'd115,  14'd538,  14'd144,  -14'd1682,  
14'd242,  -14'd300,  14'd138,  -14'd75,  14'd1435,  -14'd1617,  14'd743,  -14'd350,  -14'd423,  -14'd756,  -14'd792,  -14'd126,  -14'd592,  -14'd18,  14'd1050,  14'd590,  
14'd1760,  14'd342,  14'd1714,  14'd264,  14'd552,  -14'd1142,  14'd1041,  -14'd298,  -14'd249,  -14'd237,  14'd147,  14'd216,  14'd283,  14'd1400,  14'd1627,  -14'd74,  
14'd1220,  14'd743,  14'd924,  14'd9,  -14'd1571,  14'd966,  -14'd238,  14'd476,  -14'd361,  14'd545,  -14'd483,  -14'd407,  -14'd378,  14'd516,  14'd597,  -14'd596,  
-14'd183,  -14'd773,  14'd2037,  14'd1118,  -14'd371,  -14'd670,  14'd412,  14'd752,  -14'd673,  14'd1138,  14'd627,  -14'd1565,  -14'd217,  14'd909,  14'd1015,  -14'd735,  
14'd1392,  14'd564,  14'd2054,  14'd426,  -14'd1117,  -14'd148,  -14'd336,  14'd359,  -14'd1498,  -14'd1297,  -14'd1589,  -14'd662,  14'd539,  -14'd211,  14'd831,  -14'd259,  
14'd845,  -14'd631,  14'd792,  14'd45,  -14'd991,  14'd544,  -14'd49,  14'd299,  -14'd240,  14'd630,  14'd521,  -14'd29,  -14'd914,  -14'd685,  -14'd492,  -14'd391,  
14'd550,  14'd711,  14'd679,  14'd302,  -14'd494,  -14'd394,  14'd1576,  -14'd97,  -14'd494,  -14'd453,  14'd549,  -14'd1114,  -14'd1527,  14'd1521,  14'd1132,  14'd1389,  
-14'd419,  14'd591,  -14'd378,  -14'd1458,  -14'd752,  -14'd96,  14'd228,  -14'd42,  14'd403,  -14'd856,  -14'd770,  -14'd671,  -14'd1419,  14'd482,  14'd1716,  14'd854,  
14'd1055,  -14'd1328,  14'd582,  14'd970,  -14'd480,  -14'd386,  -14'd283,  -14'd1171,  -14'd1285,  14'd874,  -14'd1077,  14'd399,  -14'd808,  14'd311,  14'd393,  -14'd60,  
14'd34,  -14'd462,  14'd837,  14'd114,  -14'd687,  14'd1048,  14'd141,  14'd342,  14'd755,  -14'd672,  -14'd457,  14'd143,  -14'd557,  14'd293,  -14'd223,  -14'd454,  
-14'd1360,  14'd0,  -14'd33,  -14'd538,  -14'd513,  -14'd429,  14'd740,  -14'd967,  -14'd1028,  -14'd697,  14'd323,  14'd845,  -14'd605,  -14'd684,  -14'd310,  -14'd1812,  
-14'd1276,  14'd690,  14'd661,  14'd276,  -14'd704,  14'd764,  14'd762,  -14'd525,  -14'd390,  -14'd865,  -14'd675,  -14'd499,  -14'd138,  14'd1231,  14'd1032,  14'd458,  
-14'd1636,  -14'd947,  14'd906,  14'd50,  -14'd1595,  14'd1300,  14'd1052,  -14'd36,  -14'd779,  14'd214,  14'd1085,  14'd625,  14'd88,  14'd9,  14'd497,  -14'd979,  
14'd1965,  -14'd2292,  14'd2079,  14'd1020,  -14'd1001,  14'd1662,  -14'd663,  14'd20,  -14'd40,  -14'd53,  14'd2003,  -14'd933,  14'd629,  14'd183,  -14'd503,  14'd696,  
14'd1075,  -14'd519,  -14'd1584,  14'd467,  -14'd271,  -14'd369,  14'd19,  14'd1887,  -14'd664,  14'd265,  -14'd1216,  14'd355,  -14'd5,  -14'd1133,  -14'd400,  -14'd706,  

-14'd558,  -14'd236,  -14'd169,  -14'd124,  -14'd728,  -14'd470,  -14'd1535,  -14'd260,  14'd506,  14'd524,  -14'd193,  14'd146,  14'd215,  14'd1157,  14'd433,  -14'd206,  
-14'd1012,  -14'd164,  -14'd176,  14'd741,  14'd674,  14'd165,  14'd848,  14'd553,  -14'd115,  -14'd1252,  14'd762,  14'd455,  14'd594,  14'd298,  14'd1312,  -14'd287,  
-14'd788,  14'd552,  14'd127,  -14'd730,  -14'd1080,  14'd63,  14'd567,  -14'd1743,  14'd68,  14'd521,  14'd570,  14'd1155,  -14'd335,  14'd1214,  -14'd231,  -14'd260,  
14'd483,  -14'd1040,  -14'd565,  -14'd1345,  14'd1309,  -14'd278,  14'd90,  14'd799,  14'd768,  -14'd184,  -14'd758,  14'd1037,  -14'd223,  -14'd473,  14'd714,  -14'd424,  
-14'd576,  -14'd167,  -14'd551,  -14'd220,  14'd165,  14'd75,  -14'd752,  14'd400,  -14'd1100,  14'd802,  -14'd339,  -14'd796,  14'd763,  -14'd995,  14'd2,  14'd670,  
-14'd814,  -14'd427,  -14'd1093,  14'd784,  14'd416,  -14'd753,  -14'd403,  -14'd22,  14'd1222,  14'd288,  14'd490,  14'd606,  14'd860,  -14'd354,  -14'd495,  -14'd781,  
-14'd1180,  -14'd609,  14'd162,  -14'd369,  -14'd39,  -14'd962,  -14'd798,  14'd977,  14'd96,  -14'd835,  14'd77,  -14'd597,  14'd826,  14'd159,  -14'd282,  -14'd375,  
-14'd64,  -14'd693,  -14'd892,  -14'd155,  14'd206,  -14'd593,  -14'd281,  14'd294,  -14'd1331,  14'd65,  -14'd910,  -14'd646,  -14'd53,  -14'd1212,  -14'd114,  14'd636,  
-14'd719,  -14'd1183,  14'd519,  14'd767,  -14'd752,  -14'd266,  -14'd181,  -14'd771,  14'd1445,  14'd306,  -14'd275,  -14'd799,  -14'd630,  14'd214,  -14'd26,  14'd0,  
-14'd517,  -14'd601,  -14'd147,  14'd923,  -14'd680,  -14'd419,  14'd1298,  -14'd770,  14'd458,  -14'd87,  -14'd247,  -14'd1209,  14'd354,  14'd878,  -14'd318,  -14'd179,  
14'd1166,  -14'd1097,  -14'd1472,  14'd426,  -14'd662,  14'd901,  -14'd798,  -14'd1001,  14'd1059,  -14'd687,  -14'd1862,  -14'd896,  -14'd1048,  -14'd1130,  14'd933,  -14'd458,  
-14'd112,  -14'd1709,  14'd444,  14'd724,  14'd1075,  -14'd229,  14'd125,  -14'd159,  -14'd920,  14'd1134,  14'd729,  -14'd60,  -14'd163,  14'd628,  -14'd99,  -14'd270,  
14'd905,  -14'd566,  -14'd605,  -14'd315,  -14'd455,  14'd73,  -14'd1341,  -14'd832,  -14'd766,  -14'd525,  -14'd986,  14'd365,  14'd471,  14'd351,  14'd82,  -14'd194,  
-14'd635,  -14'd1213,  14'd311,  -14'd772,  -14'd824,  -14'd1513,  -14'd1511,  14'd82,  -14'd184,  -14'd667,  14'd1210,  -14'd771,  -14'd96,  -14'd735,  -14'd639,  14'd43,  
14'd467,  -14'd321,  -14'd985,  -14'd401,  14'd651,  -14'd1088,  14'd795,  14'd46,  -14'd55,  -14'd175,  -14'd313,  -14'd890,  14'd241,  -14'd324,  -14'd301,  14'd85,  
14'd849,  -14'd1066,  -14'd1014,  -14'd131,  14'd706,  -14'd717,  14'd662,  14'd389,  -14'd45,  14'd1143,  -14'd222,  -14'd361,  -14'd568,  -14'd1211,  -14'd652,  -14'd280,  
-14'd553,  -14'd298,  -14'd1422,  14'd140,  -14'd1019,  -14'd601,  -14'd750,  -14'd486,  -14'd358,  -14'd678,  -14'd502,  14'd67,  14'd153,  -14'd877,  -14'd915,  14'd921,  
14'd139,  -14'd464,  14'd482,  -14'd1245,  14'd1115,  -14'd113,  -14'd1697,  -14'd69,  -14'd99,  -14'd1598,  -14'd15,  -14'd680,  14'd930,  -14'd749,  -14'd353,  -14'd445,  
14'd93,  14'd710,  14'd987,  -14'd602,  -14'd1362,  -14'd1053,  -14'd113,  14'd287,  14'd1010,  -14'd83,  14'd677,  -14'd520,  14'd602,  14'd1210,  -14'd423,  14'd819,  
14'd43,  -14'd1324,  14'd657,  14'd536,  -14'd150,  -14'd1096,  -14'd546,  14'd1450,  -14'd1162,  -14'd1640,  -14'd969,  14'd258,  -14'd375,  -14'd1197,  14'd384,  -14'd188,  
14'd966,  -14'd390,  -14'd1030,  -14'd334,  14'd111,  14'd112,  14'd494,  -14'd518,  14'd728,  -14'd37,  14'd88,  14'd135,  14'd382,  -14'd1179,  -14'd580,  14'd72,  
14'd479,  14'd551,  -14'd681,  14'd1145,  -14'd1453,  14'd1054,  -14'd266,  -14'd952,  -14'd472,  -14'd387,  -14'd653,  -14'd694,  14'd747,  -14'd163,  14'd573,  14'd634,  
14'd29,  -14'd1664,  14'd66,  14'd302,  -14'd482,  -14'd92,  -14'd189,  14'd690,  14'd7,  -14'd624,  14'd1071,  -14'd1731,  14'd440,  14'd864,  -14'd552,  -14'd524,  
14'd672,  14'd95,  -14'd882,  -14'd403,  14'd832,  -14'd1380,  -14'd668,  -14'd551,  14'd784,  -14'd1540,  -14'd1091,  14'd661,  14'd690,  14'd279,  14'd379,  14'd975,  
-14'd1599,  -14'd388,  -14'd1499,  14'd46,  -14'd1304,  14'd359,  -14'd1421,  -14'd385,  14'd873,  -14'd653,  -14'd105,  14'd1090,  -14'd182,  -14'd751,  -14'd1490,  -14'd370,  

14'd242,  14'd469,  -14'd499,  14'd156,  14'd803,  14'd1310,  -14'd486,  -14'd686,  -14'd1268,  14'd397,  14'd1726,  -14'd840,  14'd1485,  -14'd193,  -14'd1432,  14'd14,  
-14'd391,  -14'd386,  -14'd1665,  14'd1819,  -14'd91,  -14'd1512,  -14'd2604,  14'd0,  14'd811,  14'd149,  -14'd614,  -14'd440,  14'd694,  -14'd3190,  14'd418,  14'd402,  
-14'd379,  14'd1652,  14'd1257,  14'd1850,  14'd501,  -14'd93,  -14'd1000,  -14'd659,  14'd417,  14'd1045,  14'd27,  14'd738,  -14'd1118,  -14'd1647,  14'd1631,  14'd210,  
14'd147,  14'd92,  14'd687,  -14'd521,  -14'd204,  14'd170,  14'd511,  -14'd999,  -14'd265,  14'd250,  -14'd319,  14'd1386,  14'd903,  14'd2343,  14'd372,  -14'd209,  
-14'd1741,  -14'd1261,  14'd41,  -14'd177,  14'd147,  -14'd779,  14'd267,  14'd273,  14'd1974,  -14'd330,  14'd138,  14'd1464,  -14'd1643,  -14'd835,  -14'd1236,  -14'd1003,  
14'd250,  14'd700,  -14'd1078,  14'd300,  14'd756,  -14'd773,  -14'd786,  -14'd798,  14'd316,  14'd83,  -14'd98,  -14'd428,  14'd306,  -14'd2389,  14'd649,  14'd732,  
-14'd1285,  14'd738,  -14'd1675,  -14'd801,  14'd1526,  14'd461,  14'd1010,  -14'd738,  -14'd100,  14'd1122,  -14'd235,  14'd448,  -14'd486,  -14'd2018,  -14'd229,  -14'd782,  
14'd221,  14'd886,  -14'd75,  -14'd103,  14'd804,  14'd96,  -14'd940,  14'd475,  -14'd2053,  -14'd17,  14'd51,  14'd676,  -14'd125,  14'd626,  -14'd1374,  14'd2291,  
14'd582,  -14'd53,  14'd280,  -14'd1684,  14'd630,  14'd1542,  14'd1909,  -14'd1857,  -14'd1489,  -14'd586,  -14'd224,  14'd1078,  14'd439,  14'd1650,  -14'd1130,  14'd1486,  
14'd39,  14'd98,  14'd51,  -14'd855,  14'd622,  14'd499,  14'd1340,  -14'd318,  -14'd1131,  -14'd2311,  14'd336,  -14'd991,  14'd255,  14'd1364,  14'd462,  -14'd1091,  
-14'd646,  14'd875,  -14'd1496,  -14'd189,  14'd1059,  14'd606,  -14'd629,  -14'd116,  14'd1826,  -14'd551,  14'd769,  14'd535,  -14'd1022,  -14'd807,  14'd124,  14'd811,  
-14'd399,  -14'd489,  -14'd990,  14'd523,  14'd1759,  14'd421,  -14'd603,  -14'd949,  14'd248,  14'd1041,  -14'd1397,  -14'd682,  -14'd177,  -14'd399,  14'd596,  14'd326,  
14'd577,  -14'd362,  14'd618,  -14'd168,  -14'd988,  -14'd292,  -14'd1240,  14'd570,  14'd337,  -14'd711,  -14'd511,  14'd695,  14'd1236,  -14'd336,  14'd1586,  -14'd924,  
14'd646,  14'd319,  14'd757,  14'd941,  -14'd401,  -14'd175,  14'd237,  -14'd1390,  14'd1103,  14'd104,  14'd656,  14'd1192,  14'd957,  14'd46,  -14'd541,  14'd296,  
14'd944,  -14'd327,  14'd230,  14'd1148,  14'd876,  -14'd513,  14'd747,  14'd232,  14'd154,  14'd543,  -14'd603,  14'd548,  14'd2334,  14'd351,  -14'd1260,  14'd229,  
-14'd684,  14'd296,  -14'd1696,  -14'd692,  14'd34,  -14'd377,  -14'd236,  -14'd836,  -14'd121,  14'd636,  14'd979,  14'd423,  -14'd250,  -14'd883,  14'd639,  14'd50,  
14'd302,  14'd280,  -14'd44,  -14'd284,  14'd202,  14'd247,  -14'd864,  -14'd1469,  14'd2352,  -14'd714,  14'd134,  14'd964,  14'd1504,  -14'd1278,  -14'd437,  -14'd261,  
-14'd867,  14'd1497,  14'd1008,  -14'd442,  14'd219,  14'd471,  -14'd542,  14'd561,  14'd169,  14'd1134,  -14'd36,  -14'd1161,  14'd1125,  -14'd1951,  -14'd607,  14'd1539,  
-14'd690,  -14'd1109,  -14'd1664,  14'd106,  14'd66,  14'd216,  14'd172,  14'd1054,  14'd73,  -14'd187,  14'd1639,  14'd437,  14'd1033,  -14'd1323,  -14'd432,  -14'd1097,  
-14'd546,  14'd1261,  -14'd1629,  14'd468,  14'd859,  -14'd1551,  -14'd658,  -14'd301,  14'd615,  14'd2101,  14'd485,  -14'd306,  14'd892,  -14'd298,  14'd984,  -14'd778,  
-14'd48,  -14'd1281,  -14'd489,  -14'd751,  -14'd234,  14'd992,  -14'd917,  -14'd624,  14'd998,  -14'd127,  14'd571,  14'd711,  -14'd251,  -14'd444,  14'd1754,  -14'd39,  
14'd873,  14'd838,  14'd646,  -14'd40,  14'd186,  -14'd559,  -14'd980,  14'd386,  14'd214,  -14'd848,  14'd361,  14'd578,  14'd383,  14'd330,  -14'd136,  14'd586,  
14'd270,  -14'd466,  -14'd357,  -14'd43,  14'd1272,  14'd328,  -14'd811,  -14'd618,  -14'd614,  14'd1097,  -14'd601,  14'd1364,  -14'd1516,  14'd140,  14'd315,  14'd1017,  
-14'd263,  14'd1051,  14'd624,  14'd169,  14'd1076,  14'd1485,  14'd590,  14'd606,  -14'd69,  -14'd552,  -14'd670,  14'd524,  -14'd80,  14'd719,  14'd391,  -14'd477,  
-14'd598,  -14'd784,  14'd354,  14'd828,  14'd104,  -14'd662,  14'd935,  -14'd786,  -14'd24,  14'd1798,  -14'd761,  14'd316,  14'd772,  14'd62,  -14'd1014,  14'd431,  

14'd841,  -14'd653,  14'd968,  -14'd1258,  -14'd1615,  -14'd755,  -14'd165,  14'd332,  14'd1441,  14'd841,  -14'd334,  14'd1201,  -14'd161,  -14'd100,  14'd237,  -14'd872,  
14'd839,  -14'd235,  -14'd760,  14'd704,  -14'd1003,  -14'd225,  14'd568,  14'd1293,  14'd131,  -14'd1110,  -14'd679,  14'd710,  -14'd111,  -14'd234,  -14'd744,  -14'd190,  
-14'd1370,  -14'd18,  -14'd737,  14'd374,  14'd251,  14'd436,  14'd349,  -14'd109,  -14'd1029,  14'd288,  -14'd1038,  14'd1304,  -14'd14,  14'd433,  -14'd630,  -14'd718,  
-14'd37,  14'd352,  14'd712,  -14'd1558,  -14'd78,  -14'd40,  14'd1020,  14'd522,  14'd283,  14'd1421,  -14'd503,  14'd1433,  -14'd775,  -14'd620,  14'd397,  -14'd610,  
14'd1295,  14'd107,  14'd1886,  14'd375,  -14'd1258,  14'd771,  -14'd1286,  14'd1098,  -14'd607,  14'd1082,  14'd630,  14'd641,  -14'd514,  -14'd681,  14'd980,  14'd1500,  
14'd384,  -14'd578,  -14'd57,  -14'd12,  14'd721,  -14'd49,  -14'd1010,  14'd1728,  14'd1865,  14'd1522,  -14'd1029,  14'd702,  14'd590,  14'd278,  14'd1319,  -14'd1015,  
-14'd813,  -14'd901,  -14'd77,  14'd817,  -14'd147,  14'd217,  14'd947,  14'd930,  14'd1303,  -14'd91,  14'd363,  14'd62,  14'd477,  14'd82,  14'd90,  -14'd96,  
-14'd198,  -14'd746,  14'd373,  14'd228,  -14'd958,  14'd692,  -14'd642,  14'd118,  14'd256,  14'd547,  -14'd255,  14'd678,  14'd1308,  -14'd806,  14'd115,  14'd478,  
-14'd843,  14'd1012,  14'd654,  -14'd292,  -14'd338,  -14'd700,  14'd186,  14'd581,  14'd248,  -14'd967,  -14'd545,  14'd87,  14'd673,  -14'd352,  14'd145,  14'd729,  
14'd1825,  -14'd30,  14'd986,  -14'd4,  14'd537,  -14'd1491,  -14'd1010,  14'd765,  -14'd622,  14'd221,  14'd686,  14'd372,  14'd1891,  14'd63,  -14'd240,  14'd2014,  
14'd464,  14'd1250,  14'd321,  14'd363,  14'd2325,  14'd825,  -14'd573,  14'd1581,  -14'd244,  -14'd1605,  -14'd576,  -14'd175,  14'd1672,  14'd984,  -14'd622,  14'd489,  
-14'd122,  14'd473,  14'd1389,  14'd1615,  14'd482,  -14'd277,  14'd1591,  14'd195,  14'd667,  -14'd1941,  14'd513,  -14'd771,  14'd59,  14'd249,  -14'd905,  14'd541,  
-14'd245,  14'd814,  -14'd298,  -14'd264,  -14'd197,  14'd933,  14'd218,  -14'd48,  14'd549,  -14'd1640,  14'd777,  14'd453,  -14'd9,  -14'd2167,  14'd396,  -14'd361,  
14'd759,  -14'd167,  -14'd1159,  14'd337,  -14'd811,  -14'd1631,  -14'd1046,  14'd216,  -14'd1711,  -14'd1476,  14'd1,  14'd697,  14'd943,  14'd1882,  14'd658,  -14'd1076,  
14'd1909,  -14'd145,  -14'd114,  14'd1137,  -14'd193,  14'd702,  14'd798,  -14'd703,  -14'd1014,  -14'd1073,  14'd7,  -14'd653,  14'd2028,  -14'd879,  -14'd679,  14'd1059,  
14'd208,  14'd734,  -14'd947,  -14'd752,  -14'd241,  14'd1083,  -14'd573,  -14'd362,  -14'd1276,  -14'd983,  -14'd1262,  14'd1959,  -14'd73,  -14'd169,  -14'd699,  -14'd766,  
-14'd209,  -14'd300,  -14'd523,  -14'd397,  14'd761,  -14'd958,  -14'd829,  -14'd136,  14'd140,  14'd722,  -14'd1669,  -14'd47,  -14'd202,  14'd979,  14'd429,  14'd1024,  
-14'd1511,  14'd1301,  -14'd717,  -14'd219,  14'd207,  -14'd104,  14'd169,  -14'd1532,  -14'd561,  -14'd658,  14'd686,  14'd40,  -14'd580,  -14'd588,  -14'd116,  14'd488,  
-14'd96,  -14'd556,  -14'd786,  -14'd339,  14'd94,  14'd1152,  -14'd923,  14'd140,  -14'd515,  14'd447,  14'd686,  14'd174,  14'd944,  14'd68,  14'd125,  14'd782,  
-14'd786,  -14'd237,  14'd2445,  -14'd1170,  14'd438,  -14'd386,  14'd34,  14'd513,  -14'd495,  14'd88,  14'd641,  14'd331,  14'd885,  14'd570,  -14'd915,  -14'd773,  
14'd773,  14'd1702,  14'd1177,  -14'd295,  14'd124,  -14'd248,  -14'd2502,  -14'd10,  -14'd1660,  14'd856,  -14'd460,  14'd1017,  14'd860,  14'd800,  14'd551,  -14'd1476,  
14'd21,  -14'd878,  -14'd963,  -14'd195,  -14'd192,  -14'd1372,  -14'd1925,  -14'd87,  -14'd1043,  14'd301,  -14'd1131,  -14'd8,  -14'd554,  14'd1144,  14'd703,  14'd430,  
-14'd568,  14'd119,  -14'd46,  -14'd433,  14'd271,  -14'd167,  14'd371,  14'd240,  -14'd1468,  -14'd2014,  -14'd526,  -14'd141,  -14'd581,  -14'd590,  -14'd482,  -14'd774,  
14'd1826,  -14'd742,  -14'd566,  -14'd50,  14'd10,  14'd343,  -14'd1148,  -14'd731,  -14'd93,  -14'd524,  -14'd279,  14'd1348,  14'd101,  14'd1715,  14'd457,  -14'd112,  
14'd496,  -14'd149,  14'd1024,  14'd1168,  14'd599,  -14'd27,  14'd930,  -14'd825,  -14'd447,  -14'd2451,  -14'd1421,  14'd391,  14'd672,  14'd419,  -14'd777,  -14'd500,  

-14'd1011,  14'd65,  14'd443,  14'd381,  14'd690,  14'd701,  -14'd2588,  14'd61,  -14'd136,  -14'd209,  -14'd622,  14'd978,  -14'd218,  14'd141,  14'd279,  -14'd319,  
14'd650,  -14'd369,  -14'd45,  -14'd1093,  14'd78,  -14'd4,  14'd692,  -14'd220,  14'd568,  -14'd746,  -14'd269,  -14'd229,  14'd1363,  -14'd1535,  14'd1203,  -14'd278,  
-14'd659,  14'd915,  14'd457,  14'd412,  -14'd663,  -14'd710,  -14'd237,  14'd346,  14'd566,  -14'd1663,  -14'd1386,  -14'd292,  14'd777,  14'd443,  14'd385,  14'd374,  
14'd134,  14'd2156,  14'd163,  -14'd964,  14'd830,  14'd225,  -14'd1628,  -14'd94,  14'd1359,  14'd864,  -14'd1713,  -14'd725,  14'd336,  -14'd543,  14'd1413,  14'd1142,  
14'd1358,  -14'd560,  14'd873,  14'd859,  -14'd465,  14'd54,  -14'd1639,  14'd703,  14'd493,  14'd1025,  -14'd1080,  14'd178,  -14'd794,  -14'd900,  -14'd138,  -14'd2685,  
-14'd614,  14'd1473,  14'd376,  -14'd199,  14'd608,  14'd232,  14'd1305,  -14'd821,  14'd50,  -14'd724,  14'd232,  -14'd292,  14'd772,  14'd993,  14'd294,  14'd707,  
14'd386,  -14'd330,  -14'd939,  14'd876,  14'd396,  14'd217,  14'd1915,  14'd339,  14'd56,  -14'd910,  14'd1296,  14'd193,  14'd69,  -14'd1769,  -14'd903,  14'd45,  
-14'd1395,  14'd2376,  -14'd956,  -14'd59,  14'd831,  14'd86,  14'd645,  14'd446,  -14'd172,  -14'd318,  -14'd675,  14'd430,  14'd167,  14'd277,  -14'd1670,  -14'd643,  
-14'd1134,  14'd3169,  -14'd188,  14'd858,  14'd1040,  -14'd1234,  -14'd512,  -14'd150,  14'd791,  -14'd295,  14'd19,  14'd1317,  14'd266,  -14'd483,  14'd1182,  14'd489,  
14'd1790,  14'd1812,  14'd1637,  -14'd763,  14'd1117,  14'd641,  14'd130,  -14'd1542,  -14'd676,  -14'd305,  14'd259,  14'd615,  14'd544,  -14'd500,  14'd654,  14'd502,  
14'd1160,  14'd965,  14'd815,  14'd765,  -14'd459,  14'd748,  14'd282,  14'd283,  -14'd1150,  -14'd1096,  -14'd954,  14'd1448,  14'd856,  14'd396,  -14'd268,  14'd862,  
-14'd388,  -14'd65,  -14'd448,  14'd149,  14'd688,  -14'd534,  14'd802,  14'd426,  14'd1850,  -14'd2050,  -14'd326,  -14'd543,  -14'd1072,  -14'd700,  -14'd363,  14'd240,  
-14'd915,  14'd436,  14'd626,  14'd820,  14'd1621,  -14'd1696,  14'd156,  14'd633,  -14'd629,  14'd229,  -14'd88,  14'd428,  -14'd1299,  14'd373,  -14'd206,  -14'd44,  
14'd1024,  -14'd41,  -14'd364,  14'd1055,  -14'd1542,  14'd1035,  -14'd346,  14'd560,  -14'd619,  -14'd885,  14'd370,  14'd648,  -14'd416,  14'd1278,  14'd799,  14'd776,  
14'd2349,  14'd1166,  14'd763,  -14'd72,  -14'd2183,  14'd207,  14'd1579,  14'd678,  14'd516,  -14'd225,  -14'd323,  14'd813,  -14'd451,  -14'd294,  14'd1580,  -14'd1132,  
-14'd210,  -14'd386,  -14'd83,  14'd217,  -14'd631,  -14'd397,  14'd1260,  14'd31,  -14'd1140,  -14'd1078,  -14'd224,  -14'd866,  -14'd1246,  -14'd446,  14'd96,  -14'd820,  
14'd902,  14'd20,  -14'd1564,  14'd1381,  14'd235,  14'd390,  14'd785,  -14'd676,  14'd725,  -14'd423,  -14'd1478,  -14'd117,  -14'd840,  -14'd1124,  14'd1429,  14'd147,  
14'd380,  14'd638,  -14'd717,  14'd120,  -14'd275,  14'd852,  14'd1288,  -14'd363,  14'd1362,  14'd1176,  14'd89,  -14'd746,  -14'd318,  -14'd389,  -14'd213,  -14'd1648,  
14'd1363,  14'd1306,  14'd1532,  14'd436,  -14'd160,  14'd1393,  14'd27,  14'd682,  -14'd311,  14'd718,  14'd341,  -14'd295,  14'd773,  -14'd552,  14'd459,  -14'd116,  
14'd377,  -14'd30,  -14'd372,  14'd442,  14'd179,  14'd395,  -14'd59,  14'd261,  14'd190,  -14'd586,  14'd324,  -14'd861,  14'd1325,  -14'd995,  14'd313,  14'd1478,  
14'd353,  14'd421,  14'd887,  -14'd401,  -14'd949,  -14'd1533,  -14'd1578,  -14'd697,  -14'd2017,  14'd1064,  -14'd2724,  14'd239,  -14'd597,  14'd0,  -14'd654,  -14'd1422,  
14'd956,  14'd759,  14'd1674,  14'd159,  -14'd465,  14'd1936,  -14'd44,  -14'd411,  -14'd302,  14'd950,  -14'd621,  -14'd372,  14'd80,  14'd1599,  14'd393,  14'd310,  
-14'd767,  -14'd401,  -14'd212,  14'd705,  -14'd221,  14'd171,  -14'd1012,  14'd369,  14'd170,  -14'd79,  14'd202,  -14'd566,  14'd960,  -14'd644,  14'd7,  -14'd1349,  
-14'd1610,  -14'd1038,  -14'd937,  -14'd402,  14'd1936,  14'd7,  14'd929,  14'd758,  -14'd2355,  14'd899,  -14'd1359,  -14'd183,  -14'd452,  -14'd697,  14'd1326,  14'd582,  
-14'd1749,  -14'd411,  -14'd2465,  14'd851,  14'd764,  14'd66,  -14'd387,  14'd392,  -14'd1326,  -14'd315,  -14'd213,  -14'd1034,  -14'd1093,  -14'd674,  -14'd707,  14'd74,  

-14'd957,  14'd2193,  -14'd847,  -14'd67,  14'd1238,  14'd1307,  -14'd724,  14'd682,  -14'd1735,  -14'd620,  -14'd400,  -14'd162,  14'd911,  -14'd505,  14'd293,  14'd820,  
14'd347,  14'd1854,  -14'd928,  -14'd9,  14'd1344,  14'd2104,  -14'd1833,  -14'd1092,  -14'd514,  14'd679,  -14'd414,  14'd112,  14'd68,  14'd420,  14'd1272,  14'd1955,  
-14'd56,  14'd130,  14'd738,  -14'd1058,  14'd826,  -14'd595,  14'd2089,  14'd51,  -14'd324,  -14'd840,  14'd32,  14'd845,  14'd461,  14'd1842,  -14'd960,  -14'd201,  
-14'd1019,  -14'd865,  14'd996,  -14'd112,  -14'd1735,  -14'd427,  -14'd247,  -14'd780,  14'd1259,  14'd90,  14'd950,  14'd44,  -14'd1119,  14'd1718,  -14'd899,  14'd586,  
-14'd2290,  -14'd2438,  14'd827,  -14'd123,  -14'd1333,  -14'd1431,  14'd42,  -14'd1034,  -14'd20,  -14'd776,  -14'd393,  -14'd1319,  -14'd1831,  -14'd776,  14'd404,  -14'd101,  
-14'd34,  -14'd508,  14'd428,  14'd42,  -14'd457,  -14'd454,  -14'd1139,  14'd1128,  -14'd1107,  -14'd64,  14'd691,  14'd637,  14'd977,  -14'd962,  -14'd1246,  14'd1749,  
14'd1254,  14'd2621,  -14'd1561,  -14'd112,  14'd285,  14'd361,  -14'd560,  14'd845,  14'd591,  -14'd959,  -14'd1269,  14'd362,  14'd712,  14'd896,  14'd646,  14'd928,  
14'd442,  14'd136,  -14'd433,  -14'd181,  -14'd915,  -14'd431,  14'd1755,  -14'd56,  -14'd463,  -14'd1119,  14'd732,  14'd473,  14'd599,  14'd838,  -14'd32,  14'd411,  
14'd942,  14'd166,  14'd1806,  -14'd1579,  14'd769,  -14'd219,  14'd1744,  14'd456,  14'd557,  14'd398,  14'd219,  14'd698,  -14'd1918,  14'd1686,  -14'd1361,  14'd634,  
14'd127,  -14'd55,  14'd1595,  14'd117,  -14'd463,  14'd67,  14'd998,  14'd1127,  -14'd474,  -14'd577,  -14'd894,  14'd1035,  14'd435,  -14'd1935,  -14'd1339,  -14'd1623,  
-14'd926,  14'd651,  -14'd730,  14'd373,  -14'd282,  -14'd1010,  -14'd1539,  -14'd437,  -14'd578,  -14'd677,  14'd1678,  -14'd762,  -14'd920,  14'd102,  14'd102,  14'd169,  
14'd1819,  14'd206,  -14'd454,  -14'd309,  -14'd1137,  14'd729,  -14'd1692,  -14'd11,  -14'd262,  -14'd480,  -14'd1437,  14'd1480,  -14'd636,  14'd359,  -14'd191,  -14'd984,  
-14'd116,  14'd46,  14'd1043,  -14'd988,  -14'd343,  14'd711,  14'd801,  14'd1749,  14'd954,  -14'd1416,  14'd42,  -14'd782,  -14'd368,  -14'd119,  14'd242,  14'd893,  
-14'd665,  14'd1067,  -14'd145,  14'd1476,  14'd962,  14'd158,  14'd540,  14'd145,  14'd391,  14'd636,  -14'd660,  -14'd1139,  14'd181,  -14'd18,  -14'd807,  -14'd804,  
-14'd77,  -14'd1391,  14'd764,  14'd989,  -14'd310,  -14'd55,  -14'd1835,  -14'd139,  14'd1263,  14'd715,  14'd485,  14'd1192,  -14'd438,  -14'd750,  14'd643,  14'd1242,  
14'd0,  -14'd61,  14'd1032,  14'd1052,  -14'd1343,  14'd120,  14'd542,  14'd1121,  14'd1039,  -14'd701,  14'd984,  -14'd1222,  -14'd90,  14'd539,  -14'd488,  -14'd917,  
14'd1097,  -14'd1152,  14'd787,  -14'd277,  14'd965,  14'd156,  14'd1970,  -14'd213,  -14'd513,  -14'd1520,  14'd1282,  -14'd109,  -14'd1321,  -14'd765,  14'd448,  14'd818,  
14'd15,  14'd119,  -14'd195,  -14'd1012,  -14'd217,  14'd121,  -14'd527,  14'd359,  14'd324,  -14'd734,  -14'd363,  -14'd956,  -14'd296,  -14'd163,  -14'd1422,  14'd205,  
14'd106,  -14'd627,  -14'd1964,  -14'd7,  -14'd70,  -14'd577,  -14'd2279,  14'd316,  14'd864,  14'd689,  -14'd1452,  14'd638,  -14'd192,  14'd1556,  14'd922,  14'd1770,  
14'd985,  14'd587,  14'd1206,  14'd634,  14'd787,  14'd1668,  14'd800,  -14'd381,  14'd928,  14'd2065,  14'd793,  14'd672,  14'd151,  -14'd1591,  14'd530,  14'd427,  
14'd722,  -14'd164,  14'd130,  14'd916,  -14'd431,  14'd1500,  14'd1238,  14'd428,  14'd1033,  14'd1079,  14'd943,  -14'd158,  14'd529,  -14'd327,  14'd181,  -14'd478,  
14'd732,  -14'd178,  14'd28,  14'd208,  -14'd314,  -14'd1102,  -14'd504,  -14'd154,  -14'd73,  -14'd1510,  -14'd271,  -14'd1529,  14'd780,  14'd347,  -14'd1518,  -14'd393,  
-14'd1335,  -14'd516,  -14'd686,  -14'd623,  14'd1371,  -14'd1031,  -14'd930,  -14'd28,  -14'd1480,  14'd1701,  -14'd329,  14'd923,  14'd1126,  -14'd787,  14'd258,  -14'd265,  
14'd249,  14'd605,  -14'd283,  -14'd1669,  -14'd633,  14'd198,  -14'd2365,  -14'd799,  14'd2123,  14'd1862,  -14'd831,  14'd640,  -14'd125,  -14'd932,  -14'd921,  14'd44,  
14'd947,  -14'd29,  14'd61,  -14'd424,  -14'd11,  14'd1312,  -14'd130,  -14'd21,  14'd459,  14'd364,  14'd107,  14'd962,  14'd1952,  -14'd241,  14'd1042,  -14'd171,  

-14'd1846,  -14'd2607,  -14'd1311,  -14'd1761,  14'd929,  -14'd1114,  14'd1197,  -14'd1020,  -14'd1147,  14'd1089,  -14'd1860,  -14'd211,  -14'd470,  -14'd181,  -14'd2172,  -14'd2220,  
14'd386,  14'd1032,  -14'd144,  -14'd1303,  -14'd1408,  -14'd1024,  -14'd447,  -14'd19,  -14'd2044,  -14'd685,  -14'd905,  -14'd593,  -14'd551,  14'd1962,  -14'd1262,  -14'd1039,  
14'd2458,  -14'd190,  14'd2135,  14'd1054,  -14'd973,  14'd714,  14'd1078,  -14'd409,  -14'd485,  -14'd1645,  -14'd16,  14'd25,  14'd127,  14'd1776,  -14'd1061,  -14'd1044,  
14'd685,  -14'd11,  -14'd301,  14'd568,  -14'd1207,  -14'd746,  14'd430,  14'd108,  14'd464,  -14'd189,  14'd1401,  14'd895,  -14'd727,  -14'd1404,  -14'd57,  -14'd85,  
14'd444,  14'd313,  14'd208,  14'd365,  -14'd531,  -14'd575,  -14'd133,  14'd614,  -14'd1223,  14'd801,  -14'd207,  14'd598,  14'd289,  -14'd536,  14'd555,  14'd1386,  
-14'd1850,  -14'd128,  -14'd2698,  -14'd341,  14'd147,  -14'd545,  -14'd877,  14'd46,  14'd953,  14'd250,  14'd46,  -14'd277,  -14'd50,  -14'd1357,  -14'd139,  -14'd224,  
14'd670,  14'd588,  14'd783,  14'd794,  14'd809,  -14'd422,  -14'd1733,  -14'd1470,  -14'd1461,  -14'd1246,  14'd1319,  14'd922,  -14'd163,  14'd2086,  -14'd576,  -14'd506,  
14'd1378,  -14'd23,  14'd1216,  -14'd153,  -14'd1461,  -14'd207,  -14'd794,  14'd1043,  14'd844,  14'd1108,  -14'd894,  14'd349,  -14'd1343,  14'd1004,  -14'd1103,  -14'd310,  
-14'd140,  14'd850,  14'd85,  -14'd713,  14'd466,  14'd454,  14'd576,  14'd231,  -14'd643,  14'd516,  14'd1092,  -14'd349,  14'd478,  14'd1393,  14'd1030,  -14'd49,  
-14'd12,  -14'd1665,  -14'd2222,  14'd551,  -14'd432,  -14'd1884,  14'd479,  -14'd259,  14'd1334,  -14'd1290,  -14'd74,  -14'd150,  -14'd2484,  14'd456,  14'd277,  14'd144,  
-14'd390,  14'd103,  -14'd1522,  14'd1001,  14'd486,  -14'd1041,  -14'd2844,  14'd338,  14'd776,  -14'd216,  14'd963,  -14'd317,  -14'd550,  -14'd1909,  14'd966,  14'd61,  
-14'd125,  -14'd767,  -14'd49,  -14'd550,  -14'd1590,  -14'd2469,  -14'd257,  -14'd2225,  -14'd784,  14'd763,  -14'd598,  -14'd1052,  -14'd140,  14'd1796,  -14'd653,  -14'd394,  
14'd1058,  -14'd23,  14'd865,  -14'd494,  -14'd435,  -14'd979,  14'd820,  14'd1230,  -14'd160,  -14'd212,  -14'd1158,  14'd387,  14'd722,  14'd1240,  -14'd482,  -14'd36,  
-14'd129,  14'd1174,  14'd2224,  -14'd803,  -14'd1348,  14'd769,  14'd1904,  -14'd574,  14'd1104,  -14'd1500,  -14'd25,  -14'd8,  -14'd1114,  14'd364,  -14'd171,  14'd207,  
14'd1570,  14'd1229,  -14'd1199,  14'd447,  -14'd891,  -14'd1787,  14'd656,  14'd1393,  -14'd125,  -14'd2776,  14'd1078,  -14'd630,  -14'd813,  -14'd1349,  14'd962,  -14'd2470,  
-14'd92,  14'd447,  -14'd325,  -14'd259,  14'd1388,  14'd286,  -14'd258,  14'd140,  -14'd686,  14'd788,  14'd80,  -14'd3010,  -14'd1288,  -14'd841,  -14'd508,  -14'd902,  
-14'd77,  -14'd2366,  -14'd119,  -14'd943,  14'd765,  -14'd1239,  14'd1118,  -14'd1072,  -14'd3441,  14'd1046,  14'd324,  14'd166,  14'd1111,  14'd120,  14'd1212,  -14'd748,  
-14'd25,  -14'd1332,  14'd1428,  -14'd890,  -14'd2591,  -14'd903,  14'd834,  -14'd1094,  14'd653,  -14'd776,  -14'd2669,  -14'd628,  -14'd521,  14'd1528,  -14'd218,  -14'd2905,  
14'd209,  14'd208,  14'd2344,  14'd1212,  -14'd2510,  -14'd1418,  -14'd602,  14'd88,  -14'd100,  14'd1248,  -14'd324,  14'd36,  -14'd1528,  -14'd769,  14'd489,  -14'd3205,  
14'd318,  14'd647,  -14'd182,  14'd153,  -14'd3198,  -14'd1950,  -14'd335,  -14'd96,  -14'd1794,  14'd1199,  -14'd1950,  14'd1044,  -14'd259,  -14'd257,  -14'd1146,  -14'd1966,  
14'd219,  14'd9,  -14'd838,  14'd1494,  -14'd662,  -14'd100,  14'd404,  14'd1193,  14'd284,  -14'd225,  -14'd750,  -14'd957,  -14'd428,  -14'd1044,  14'd20,  14'd772,  
14'd1635,  14'd34,  14'd688,  14'd1054,  -14'd3173,  14'd1160,  -14'd676,  -14'd80,  14'd1527,  14'd1900,  -14'd939,  -14'd221,  -14'd571,  -14'd458,  14'd2,  14'd446,  
14'd154,  -14'd821,  14'd386,  14'd490,  14'd795,  -14'd266,  14'd984,  -14'd167,  14'd1436,  14'd2598,  14'd416,  -14'd49,  -14'd596,  -14'd975,  14'd623,  14'd735,  
-14'd1145,  -14'd1375,  14'd818,  14'd959,  14'd207,  -14'd1669,  -14'd1047,  14'd816,  14'd897,  14'd158,  14'd814,  -14'd346,  -14'd134,  14'd455,  14'd629,  14'd1806,  
-14'd343,  -14'd1124,  -14'd191,  14'd504,  -14'd52,  -14'd1840,  14'd219,  14'd178,  -14'd1883,  14'd1070,  14'd380,  14'd1476,  14'd443,  14'd163,  14'd361,  14'd1490,  

14'd587,  -14'd332,  -14'd742,  -14'd22,  14'd1755,  -14'd1159,  14'd1044,  -14'd563,  -14'd218,  14'd1120,  14'd330,  -14'd100,  -14'd1306,  -14'd1159,  -14'd561,  14'd850,  
-14'd561,  -14'd144,  -14'd1777,  -14'd1189,  14'd771,  14'd397,  14'd1365,  14'd392,  14'd91,  -14'd438,  -14'd2263,  -14'd190,  14'd1385,  14'd343,  -14'd145,  -14'd157,  
-14'd37,  -14'd58,  -14'd631,  -14'd1394,  -14'd344,  -14'd39,  -14'd300,  14'd0,  -14'd755,  -14'd1325,  -14'd1260,  14'd1108,  14'd145,  14'd735,  14'd613,  14'd635,  
14'd631,  14'd688,  -14'd1242,  -14'd692,  -14'd6,  -14'd29,  14'd1037,  -14'd619,  14'd1285,  -14'd451,  -14'd77,  14'd273,  14'd508,  14'd3011,  14'd755,  14'd966,  
-14'd391,  -14'd233,  14'd116,  -14'd407,  14'd270,  14'd482,  14'd219,  14'd704,  -14'd205,  -14'd16,  14'd52,  -14'd738,  -14'd966,  14'd503,  14'd1731,  14'd522,  
14'd57,  14'd1648,  -14'd615,  -14'd949,  -14'd914,  -14'd502,  14'd1387,  -14'd1529,  -14'd613,  14'd960,  14'd1019,  14'd312,  14'd19,  -14'd2067,  -14'd17,  -14'd376,  
14'd946,  14'd967,  -14'd473,  -14'd473,  14'd171,  -14'd311,  -14'd470,  -14'd1020,  14'd931,  14'd1396,  -14'd293,  -14'd771,  -14'd632,  -14'd872,  -14'd80,  14'd229,  
-14'd172,  14'd1243,  14'd92,  -14'd1107,  14'd520,  14'd1367,  -14'd494,  14'd151,  14'd310,  -14'd293,  14'd479,  -14'd164,  -14'd59,  -14'd85,  -14'd537,  -14'd269,  
14'd890,  14'd2,  14'd1338,  14'd727,  14'd549,  14'd478,  14'd990,  14'd102,  -14'd684,  -14'd1323,  14'd120,  14'd779,  -14'd327,  14'd313,  -14'd489,  -14'd988,  
14'd40,  14'd900,  14'd1262,  14'd1217,  -14'd471,  14'd1544,  -14'd483,  14'd11,  14'd848,  -14'd578,  14'd303,  -14'd257,  -14'd1028,  14'd1079,  14'd1498,  -14'd1463,  
14'd13,  14'd703,  -14'd895,  14'd109,  -14'd1370,  14'd471,  14'd795,  -14'd268,  -14'd181,  14'd383,  -14'd1188,  14'd1956,  14'd482,  -14'd137,  14'd613,  14'd63,  
-14'd157,  -14'd89,  -14'd1018,  -14'd459,  -14'd152,  -14'd799,  -14'd288,  14'd95,  14'd2162,  14'd224,  -14'd1582,  14'd224,  -14'd1225,  -14'd15,  -14'd82,  -14'd930,  
14'd413,  14'd766,  -14'd1547,  14'd1244,  14'd991,  -14'd1104,  14'd558,  14'd97,  14'd293,  14'd55,  -14'd200,  14'd422,  -14'd538,  -14'd121,  -14'd583,  14'd800,  
14'd1388,  -14'd122,  14'd623,  14'd360,  -14'd1111,  14'd654,  14'd85,  14'd880,  14'd578,  14'd902,  -14'd131,  -14'd158,  -14'd444,  14'd507,  14'd1443,  14'd309,  
14'd912,  14'd447,  -14'd236,  14'd587,  -14'd196,  14'd1234,  14'd577,  14'd873,  -14'd404,  -14'd447,  -14'd438,  14'd94,  14'd1338,  14'd197,  14'd437,  14'd645,  
14'd924,  14'd852,  14'd1138,  14'd1620,  14'd435,  14'd231,  14'd933,  14'd986,  -14'd692,  14'd641,  14'd200,  -14'd712,  14'd662,  14'd1058,  14'd1217,  -14'd192,  
14'd1157,  -14'd423,  14'd1234,  14'd322,  -14'd926,  -14'd428,  -14'd254,  14'd230,  -14'd7,  -14'd1383,  -14'd349,  -14'd680,  -14'd759,  14'd269,  14'd914,  -14'd1151,  
14'd1213,  14'd639,  -14'd2179,  14'd630,  14'd812,  14'd225,  -14'd1122,  14'd1133,  -14'd1901,  -14'd258,  14'd853,  -14'd341,  14'd1377,  -14'd322,  -14'd3,  14'd894,  
14'd315,  -14'd1147,  14'd174,  -14'd51,  14'd1256,  14'd425,  -14'd1161,  14'd1269,  -14'd1162,  14'd115,  -14'd1161,  -14'd650,  14'd342,  14'd1266,  -14'd454,  14'd1810,  
14'd456,  14'd568,  -14'd55,  14'd1663,  14'd353,  14'd967,  14'd928,  14'd309,  14'd425,  14'd827,  14'd505,  14'd188,  14'd1120,  14'd916,  -14'd1,  -14'd499,  
14'd732,  -14'd209,  14'd663,  14'd1908,  14'd2457,  14'd1261,  -14'd1406,  14'd1358,  -14'd1491,  14'd418,  14'd97,  14'd165,  14'd1523,  14'd251,  14'd1621,  14'd129,  
-14'd1669,  14'd191,  14'd608,  14'd1544,  14'd614,  -14'd119,  -14'd565,  14'd684,  -14'd52,  -14'd250,  -14'd413,  -14'd335,  -14'd523,  14'd1511,  14'd794,  -14'd361,  
-14'd949,  14'd1253,  -14'd1104,  -14'd1115,  -14'd626,  -14'd112,  -14'd1386,  14'd557,  -14'd2267,  -14'd694,  14'd1210,  -14'd48,  -14'd316,  -14'd2134,  -14'd1254,  -14'd387,  
14'd489,  -14'd232,  14'd522,  14'd1156,  -14'd484,  14'd1027,  14'd307,  14'd1429,  14'd358,  14'd423,  -14'd618,  14'd886,  -14'd348,  -14'd928,  -14'd1454,  -14'd956,  
14'd259,  14'd8,  14'd443,  14'd510,  -14'd783,  14'd808,  14'd688,  14'd294,  14'd1581,  14'd58,  14'd139,  14'd169,  14'd1239,  -14'd975,  -14'd330,  -14'd207,  

14'd156,  14'd813,  -14'd690,  -14'd1555,  14'd124,  -14'd1080,  14'd970,  -14'd1936,  -14'd1451,  -14'd1007,  -14'd780,  14'd1175,  -14'd432,  14'd289,  -14'd135,  -14'd1398,  
14'd632,  -14'd458,  -14'd256,  -14'd700,  -14'd96,  -14'd19,  14'd98,  -14'd922,  -14'd1524,  14'd23,  -14'd315,  14'd134,  -14'd755,  14'd546,  14'd450,  14'd1205,  
14'd899,  14'd1813,  -14'd888,  -14'd420,  14'd763,  -14'd405,  14'd921,  -14'd1120,  -14'd254,  14'd969,  14'd629,  14'd840,  -14'd1451,  14'd269,  -14'd45,  14'd403,  
14'd1400,  -14'd888,  14'd912,  14'd582,  -14'd878,  -14'd707,  14'd695,  -14'd2055,  -14'd497,  14'd1292,  14'd590,  -14'd303,  -14'd194,  -14'd189,  14'd844,  14'd492,  
-14'd1179,  -14'd2676,  -14'd1006,  -14'd1334,  -14'd187,  14'd113,  14'd745,  14'd252,  -14'd1128,  -14'd1371,  -14'd572,  14'd612,  14'd311,  -14'd1331,  -14'd1127,  14'd875,  
-14'd48,  -14'd420,  14'd520,  -14'd1717,  -14'd1492,  -14'd505,  14'd365,  -14'd1338,  14'd1032,  -14'd754,  14'd1609,  14'd55,  -14'd1845,  14'd299,  -14'd753,  14'd388,  
-14'd269,  14'd969,  -14'd176,  -14'd228,  14'd543,  14'd936,  14'd99,  -14'd836,  -14'd1332,  -14'd219,  -14'd1058,  14'd236,  -14'd22,  14'd230,  -14'd1323,  -14'd1477,  
14'd432,  -14'd73,  -14'd731,  14'd495,  -14'd978,  14'd156,  14'd790,  -14'd1667,  -14'd400,  -14'd18,  -14'd762,  14'd846,  -14'd861,  -14'd113,  14'd25,  14'd1391,  
14'd901,  14'd1306,  14'd526,  -14'd2072,  -14'd811,  14'd343,  14'd1652,  14'd636,  -14'd562,  14'd1784,  14'd56,  14'd333,  14'd438,  14'd1599,  -14'd592,  14'd258,  
14'd728,  14'd1186,  14'd2112,  -14'd1166,  -14'd968,  -14'd1296,  14'd352,  -14'd864,  14'd1190,  -14'd1267,  -14'd260,  -14'd1152,  -14'd1504,  14'd67,  -14'd1087,  14'd621,  
-14'd1538,  -14'd1058,  14'd1453,  14'd815,  -14'd91,  -14'd101,  -14'd411,  14'd589,  14'd760,  14'd911,  -14'd1410,  -14'd724,  -14'd1034,  -14'd436,  14'd603,  -14'd629,  
14'd83,  14'd438,  -14'd415,  -14'd20,  -14'd1300,  14'd311,  14'd933,  14'd517,  -14'd295,  -14'd256,  14'd258,  -14'd785,  14'd482,  -14'd32,  -14'd466,  14'd39,  
14'd1482,  14'd362,  14'd2302,  -14'd161,  -14'd1506,  14'd1461,  14'd1124,  14'd634,  -14'd685,  -14'd184,  14'd363,  14'd719,  14'd489,  14'd1899,  14'd455,  14'd1223,  
14'd1191,  14'd1548,  14'd1784,  -14'd203,  -14'd1375,  -14'd643,  14'd1655,  14'd2023,  14'd843,  14'd446,  14'd924,  14'd1140,  -14'd342,  14'd1544,  14'd433,  -14'd1241,  
14'd458,  14'd468,  -14'd799,  -14'd621,  14'd166,  -14'd1098,  14'd548,  -14'd78,  -14'd970,  -14'd1481,  -14'd887,  -14'd576,  14'd510,  14'd516,  -14'd1356,  -14'd684,  
14'd969,  -14'd1400,  -14'd632,  -14'd1077,  -14'd1559,  14'd754,  14'd1159,  -14'd403,  14'd1508,  -14'd90,  14'd1241,  -14'd123,  -14'd317,  14'd535,  -14'd362,  -14'd655,  
14'd238,  14'd669,  14'd280,  14'd571,  -14'd385,  -14'd422,  14'd1373,  14'd895,  -14'd916,  -14'd818,  14'd2104,  -14'd2,  14'd957,  14'd1789,  14'd329,  14'd31,  
-14'd1414,  14'd822,  14'd1851,  -14'd348,  -14'd797,  14'd397,  14'd1611,  14'd456,  14'd634,  14'd705,  -14'd1214,  -14'd1201,  14'd730,  14'd2501,  -14'd593,  -14'd127,  
-14'd259,  -14'd1038,  14'd388,  14'd161,  14'd90,  -14'd1854,  -14'd464,  -14'd20,  -14'd1777,  -14'd1620,  -14'd1632,  -14'd65,  -14'd629,  14'd563,  -14'd1022,  -14'd693,  
14'd158,  14'd29,  14'd1195,  14'd1114,  -14'd2403,  -14'd1723,  -14'd1535,  -14'd850,  -14'd232,  -14'd373,  -14'd982,  -14'd656,  -14'd140,  14'd1595,  -14'd328,  -14'd1675,  
-14'd1245,  14'd910,  -14'd914,  -14'd1321,  14'd638,  -14'd135,  14'd2266,  14'd1029,  -14'd598,  14'd804,  14'd291,  14'd1220,  -14'd551,  -14'd2190,  -14'd508,  14'd419,  
-14'd659,  14'd280,  -14'd490,  14'd452,  14'd1244,  -14'd1133,  14'd1031,  -14'd163,  14'd1302,  14'd827,  14'd694,  -14'd1557,  -14'd793,  14'd1158,  -14'd786,  -14'd1311,  
-14'd268,  -14'd306,  14'd1267,  14'd22,  14'd903,  -14'd123,  14'd1332,  14'd1086,  14'd1572,  14'd1539,  -14'd88,  -14'd2440,  -14'd629,  14'd1338,  14'd687,  -14'd1050,  
-14'd2050,  -14'd426,  -14'd761,  14'd255,  14'd1241,  -14'd736,  -14'd965,  -14'd1258,  14'd540,  14'd1185,  14'd425,  -14'd584,  14'd253,  14'd802,  14'd189,  -14'd927,  
14'd162,  -14'd748,  14'd3382,  14'd335,  14'd1120,  14'd173,  -14'd797,  -14'd1795,  -14'd950,  14'd4971,  14'd357,  14'd2504,  14'd2227,  -14'd2304,  14'd2008,  -14'd740,  

-14'd18,  -14'd241,  14'd1379,  14'd619,  14'd417,  14'd646,  -14'd1248,  14'd1160,  14'd1364,  14'd684,  -14'd551,  14'd1727,  -14'd796,  14'd437,  -14'd125,  -14'd62,  
-14'd490,  -14'd704,  14'd1260,  14'd30,  -14'd327,  -14'd481,  -14'd1125,  14'd1222,  14'd506,  14'd508,  -14'd1093,  -14'd781,  14'd469,  14'd1156,  14'd974,  -14'd223,  
14'd1065,  -14'd2072,  14'd750,  -14'd402,  -14'd243,  -14'd286,  14'd681,  -14'd70,  14'd899,  -14'd52,  -14'd159,  -14'd791,  -14'd796,  14'd2149,  -14'd552,  -14'd405,  
-14'd1318,  -14'd1786,  -14'd1169,  -14'd1165,  -14'd690,  14'd1007,  14'd1365,  14'd404,  -14'd122,  14'd469,  14'd158,  -14'd465,  -14'd266,  14'd2268,  -14'd722,  -14'd874,  
14'd2261,  14'd2014,  -14'd250,  -14'd374,  14'd1249,  14'd441,  14'd631,  -14'd163,  14'd990,  14'd530,  14'd50,  14'd343,  -14'd548,  -14'd74,  -14'd903,  14'd44,  
-14'd895,  -14'd257,  -14'd122,  14'd1339,  14'd2481,  14'd951,  -14'd1465,  14'd792,  -14'd3,  -14'd40,  14'd64,  14'd562,  14'd795,  14'd1977,  -14'd475,  14'd1686,  
-14'd1770,  14'd1528,  14'd439,  14'd265,  -14'd1037,  -14'd1026,  14'd694,  -14'd175,  -14'd755,  -14'd51,  -14'd1346,  14'd261,  14'd616,  -14'd220,  14'd1539,  14'd359,  
14'd458,  -14'd496,  14'd402,  14'd652,  -14'd237,  -14'd29,  14'd244,  -14'd66,  14'd103,  -14'd997,  14'd1401,  -14'd11,  -14'd731,  14'd326,  -14'd51,  14'd63,  
14'd1500,  -14'd786,  14'd855,  14'd753,  -14'd216,  -14'd501,  14'd1609,  14'd1240,  14'd269,  -14'd276,  14'd17,  -14'd206,  14'd1154,  14'd419,  -14'd789,  -14'd1014,  
14'd2772,  -14'd113,  -14'd1649,  -14'd3,  -14'd1009,  -14'd644,  14'd124,  -14'd121,  -14'd227,  -14'd1511,  14'd406,  -14'd730,  14'd622,  -14'd232,  -14'd889,  14'd820,  
-14'd808,  14'd1461,  -14'd1738,  -14'd729,  -14'd404,  -14'd184,  -14'd807,  14'd928,  -14'd563,  14'd993,  14'd1034,  -14'd3,  14'd1043,  14'd308,  14'd148,  14'd30,  
-14'd268,  14'd925,  14'd323,  14'd181,  -14'd583,  14'd423,  14'd449,  -14'd667,  -14'd944,  -14'd1268,  14'd779,  -14'd99,  14'd1379,  14'd63,  14'd512,  14'd1483,  
-14'd629,  -14'd1072,  14'd606,  14'd392,  -14'd62,  14'd386,  14'd878,  14'd1203,  -14'd371,  -14'd583,  14'd204,  14'd431,  14'd1933,  -14'd597,  14'd691,  -14'd104,  
14'd687,  14'd16,  14'd821,  14'd1201,  14'd344,  -14'd1017,  14'd1164,  14'd771,  14'd135,  14'd360,  14'd1100,  -14'd304,  14'd782,  -14'd1848,  -14'd692,  -14'd922,  
-14'd1783,  -14'd570,  -14'd1331,  -14'd1328,  14'd623,  -14'd163,  14'd542,  14'd4,  -14'd1799,  14'd287,  14'd990,  -14'd481,  14'd229,  -14'd1366,  -14'd560,  14'd207,  
-14'd164,  14'd536,  -14'd1107,  -14'd830,  14'd1829,  14'd178,  -14'd506,  14'd369,  14'd727,  14'd328,  14'd1901,  14'd344,  -14'd1516,  -14'd260,  -14'd1289,  -14'd259,  
-14'd419,  14'd874,  -14'd201,  -14'd1399,  14'd764,  -14'd155,  14'd2412,  -14'd213,  -14'd268,  14'd656,  14'd581,  -14'd293,  14'd409,  -14'd809,  -14'd169,  14'd902,  
-14'd17,  14'd455,  14'd282,  14'd153,  -14'd1240,  14'd835,  14'd543,  -14'd281,  14'd1478,  14'd639,  -14'd974,  -14'd1629,  -14'd42,  14'd341,  -14'd493,  14'd174,  
14'd281,  -14'd941,  14'd229,  14'd631,  -14'd1709,  14'd790,  -14'd46,  -14'd248,  14'd218,  14'd584,  14'd1875,  14'd108,  -14'd546,  14'd1346,  -14'd157,  14'd481,  
-14'd437,  -14'd1453,  14'd691,  -14'd115,  14'd638,  14'd81,  14'd146,  14'd223,  14'd467,  -14'd1183,  14'd202,  14'd655,  -14'd430,  -14'd195,  -14'd759,  14'd495,  
-14'd1020,  -14'd1364,  -14'd1148,  14'd514,  14'd348,  -14'd178,  -14'd257,  -14'd549,  14'd1199,  14'd210,  -14'd125,  -14'd427,  14'd406,  -14'd1656,  14'd109,  -14'd80,  
-14'd812,  -14'd257,  -14'd501,  -14'd610,  -14'd861,  -14'd549,  14'd1110,  14'd1070,  14'd2158,  14'd718,  14'd769,  14'd250,  14'd155,  14'd1528,  -14'd650,  14'd1373,  
14'd1688,  14'd264,  14'd724,  14'd940,  14'd366,  -14'd767,  14'd1612,  -14'd519,  14'd225,  14'd2055,  -14'd301,  14'd231,  -14'd598,  14'd2396,  14'd279,  14'd159,  
14'd1340,  14'd327,  14'd588,  -14'd598,  14'd10,  14'd441,  -14'd143,  -14'd541,  -14'd841,  -14'd148,  14'd885,  -14'd301,  -14'd467,  14'd756,  14'd178,  14'd373,  
14'd1523,  -14'd321,  14'd745,  14'd1119,  -14'd69,  14'd44,  14'd688,  14'd312,  -14'd2014,  -14'd2308,  14'd698,  -14'd460,  -14'd140,  14'd804,  -14'd332,  14'd456,  

14'd1338,  14'd272,  14'd800,  -14'd91,  14'd240,  -14'd261,  -14'd1360,  14'd26,  14'd558,  14'd1052,  -14'd1979,  14'd362,  -14'd528,  -14'd1497,  14'd1209,  14'd1989,  
-14'd127,  14'd558,  14'd2494,  14'd237,  14'd400,  -14'd954,  14'd817,  14'd1752,  -14'd2168,  14'd457,  -14'd1777,  -14'd31,  -14'd2758,  14'd1614,  -14'd1230,  14'd8,  
-14'd732,  -14'd1922,  14'd1265,  -14'd1142,  -14'd1750,  -14'd776,  14'd1678,  14'd655,  14'd144,  14'd66,  -14'd1802,  -14'd307,  -14'd1113,  14'd1991,  14'd326,  -14'd2321,  
-14'd2006,  14'd1379,  14'd721,  -14'd835,  -14'd2013,  -14'd516,  14'd892,  -14'd119,  14'd272,  14'd262,  -14'd34,  -14'd1108,  -14'd1420,  -14'd723,  -14'd1313,  -14'd2703,  
-14'd1395,  14'd222,  -14'd830,  -14'd964,  -14'd2037,  -14'd1567,  -14'd1775,  -14'd1365,  -14'd1602,  -14'd538,  -14'd910,  -14'd1244,  -14'd2523,  -14'd1876,  14'd330,  -14'd1241,  
-14'd841,  -14'd624,  -14'd1613,  14'd1035,  14'd860,  14'd1572,  14'd1081,  -14'd564,  -14'd660,  -14'd563,  -14'd424,  14'd663,  14'd859,  -14'd83,  -14'd1508,  -14'd30,  
14'd777,  14'd1138,  14'd3249,  14'd122,  14'd0,  14'd1919,  14'd2261,  14'd1838,  -14'd860,  14'd313,  -14'd363,  14'd1064,  14'd328,  14'd1610,  14'd379,  -14'd85,  
-14'd2606,  14'd1472,  14'd259,  14'd225,  -14'd970,  14'd1181,  14'd2004,  14'd2303,  14'd339,  14'd1582,  -14'd357,  -14'd1500,  14'd1006,  -14'd275,  -14'd258,  -14'd2384,  
14'd1405,  -14'd1530,  14'd1309,  -14'd82,  -14'd277,  -14'd1259,  -14'd1897,  -14'd492,  -14'd364,  14'd1763,  -14'd1033,  14'd915,  14'd596,  14'd43,  14'd528,  14'd309,  
14'd1270,  14'd109,  14'd276,  -14'd542,  14'd725,  14'd812,  -14'd911,  -14'd1253,  14'd96,  14'd1605,  -14'd2108,  14'd1379,  -14'd1597,  -14'd1337,  14'd241,  -14'd506,  
-14'd832,  14'd358,  -14'd104,  14'd203,  14'd1008,  14'd1097,  14'd1019,  -14'd1208,  14'd42,  14'd348,  14'd124,  14'd678,  14'd207,  14'd1114,  14'd793,  14'd1286,  
-14'd1405,  14'd75,  -14'd332,  -14'd1751,  14'd802,  -14'd110,  14'd2942,  -14'd567,  -14'd1003,  -14'd471,  -14'd593,  -14'd713,  -14'd365,  14'd768,  14'd1275,  -14'd1154,  
-14'd681,  14'd1020,  14'd462,  14'd1580,  14'd391,  -14'd166,  -14'd405,  -14'd1142,  14'd810,  -14'd1222,  14'd1646,  -14'd276,  14'd393,  14'd492,  14'd210,  14'd1036,  
14'd463,  14'd735,  14'd1241,  -14'd6,  14'd77,  -14'd845,  -14'd880,  -14'd728,  14'd71,  14'd660,  14'd1022,  -14'd1183,  14'd611,  14'd1083,  14'd1355,  -14'd125,  
14'd299,  -14'd860,  14'd547,  14'd1207,  14'd433,  -14'd751,  14'd885,  -14'd906,  14'd199,  -14'd310,  14'd379,  14'd91,  14'd994,  -14'd1694,  14'd676,  14'd344,  
-14'd605,  -14'd100,  14'd967,  -14'd912,  -14'd701,  14'd332,  14'd1266,  14'd724,  14'd372,  -14'd474,  14'd1101,  -14'd732,  -14'd477,  -14'd593,  14'd205,  -14'd1373,  
-14'd894,  -14'd4,  14'd99,  -14'd620,  14'd1428,  14'd161,  14'd338,  -14'd890,  -14'd1111,  14'd328,  -14'd1361,  14'd905,  -14'd624,  -14'd268,  14'd251,  14'd682,  
14'd493,  -14'd72,  14'd1092,  -14'd1629,  14'd887,  14'd1,  14'd405,  -14'd524,  14'd653,  -14'd60,  -14'd1681,  14'd315,  -14'd1667,  14'd1622,  14'd1827,  14'd183,  
14'd2301,  -14'd1000,  14'd1295,  -14'd670,  -14'd1373,  -14'd953,  -14'd209,  -14'd1247,  14'd998,  14'd844,  14'd214,  14'd868,  -14'd54,  14'd425,  14'd914,  14'd651,  
14'd352,  14'd1628,  14'd2277,  14'd633,  -14'd7,  14'd2001,  14'd665,  -14'd495,  14'd1690,  14'd326,  -14'd810,  14'd335,  14'd435,  14'd346,  -14'd259,  -14'd379,  
14'd559,  -14'd1080,  14'd734,  -14'd2997,  -14'd802,  -14'd1698,  -14'd173,  -14'd251,  -14'd2021,  -14'd55,  -14'd1569,  -14'd767,  -14'd1365,  -14'd80,  -14'd596,  -14'd1493,  
-14'd164,  14'd223,  -14'd1333,  -14'd1256,  -14'd420,  -14'd779,  -14'd813,  -14'd979,  -14'd814,  -14'd529,  -14'd2120,  -14'd193,  -14'd1472,  -14'd956,  -14'd282,  -14'd1678,  
14'd1693,  -14'd662,  14'd694,  -14'd1506,  -14'd1914,  14'd1675,  14'd70,  14'd598,  -14'd690,  -14'd1098,  -14'd851,  -14'd1194,  14'd357,  14'd1271,  14'd813,  14'd296,  
14'd727,  14'd546,  14'd653,  -14'd108,  -14'd530,  -14'd15,  14'd634,  14'd1504,  -14'd1162,  -14'd274,  -14'd843,  -14'd645,  -14'd879,  14'd153,  14'd1943,  -14'd523,  
-14'd647,  14'd699,  14'd515,  -14'd827,  14'd984,  14'd749,  14'd951,  14'd2585,  -14'd474,  14'd76,  -14'd1317,  -14'd1296,  14'd13,  14'd1222,  -14'd97,  14'd809,  

14'd23,  14'd310,  14'd483,  -14'd518,  -14'd1353,  -14'd607,  -14'd971,  14'd202,  -14'd1530,  14'd885,  -14'd175,  14'd1256,  14'd862,  14'd627,  -14'd108,  -14'd308,  
-14'd588,  -14'd119,  -14'd1255,  -14'd607,  14'd645,  14'd1167,  -14'd407,  -14'd251,  -14'd664,  -14'd1175,  14'd1411,  14'd739,  -14'd1004,  -14'd1319,  -14'd1571,  14'd655,  
-14'd40,  -14'd473,  -14'd599,  14'd1219,  -14'd1079,  -14'd523,  14'd352,  14'd1152,  14'd47,  14'd404,  -14'd62,  -14'd118,  -14'd6,  14'd383,  14'd1320,  -14'd212,  
-14'd107,  -14'd589,  14'd474,  -14'd1411,  14'd156,  14'd853,  -14'd604,  14'd324,  -14'd334,  -14'd734,  14'd960,  14'd49,  14'd424,  -14'd1438,  14'd591,  -14'd1282,  
-14'd359,  -14'd546,  -14'd1409,  -14'd1302,  -14'd7,  -14'd564,  14'd607,  14'd324,  -14'd626,  -14'd1827,  14'd477,  14'd205,  -14'd943,  -14'd1263,  14'd740,  -14'd527,  
-14'd304,  -14'd810,  14'd287,  14'd945,  -14'd506,  -14'd190,  -14'd627,  -14'd1150,  -14'd244,  -14'd714,  -14'd1358,  -14'd345,  14'd542,  -14'd675,  14'd88,  14'd103,  
14'd370,  14'd1346,  14'd605,  -14'd949,  -14'd972,  14'd1197,  14'd90,  -14'd390,  -14'd1086,  14'd993,  -14'd549,  -14'd302,  -14'd1198,  14'd1064,  14'd84,  14'd390,  
14'd942,  14'd904,  -14'd1396,  14'd40,  14'd293,  -14'd369,  -14'd573,  -14'd556,  -14'd471,  14'd260,  -14'd1193,  -14'd1110,  -14'd33,  -14'd1109,  -14'd952,  14'd952,  
14'd112,  14'd524,  14'd472,  -14'd1282,  -14'd529,  -14'd421,  14'd895,  -14'd453,  14'd986,  -14'd1802,  -14'd223,  -14'd319,  14'd43,  -14'd486,  -14'd126,  -14'd1639,  
-14'd196,  -14'd4,  14'd1505,  14'd265,  -14'd377,  -14'd1100,  -14'd785,  -14'd556,  -14'd131,  14'd64,  -14'd467,  14'd676,  14'd97,  14'd631,  14'd826,  14'd536,  
14'd507,  14'd567,  14'd1061,  14'd260,  14'd125,  -14'd473,  14'd584,  14'd777,  -14'd1202,  -14'd842,  14'd434,  14'd1084,  -14'd1362,  -14'd1502,  14'd579,  -14'd1230,  
14'd641,  14'd252,  -14'd633,  -14'd1067,  -14'd595,  14'd897,  -14'd627,  -14'd803,  -14'd88,  14'd447,  -14'd121,  14'd404,  14'd738,  -14'd1639,  -14'd277,  -14'd415,  
-14'd718,  14'd458,  -14'd507,  -14'd395,  14'd218,  -14'd662,  14'd231,  -14'd773,  14'd124,  -14'd679,  -14'd892,  -14'd1389,  -14'd1483,  14'd685,  -14'd77,  14'd224,  
-14'd343,  -14'd1505,  -14'd171,  -14'd531,  -14'd837,  -14'd964,  -14'd243,  -14'd164,  -14'd83,  -14'd431,  14'd115,  14'd93,  14'd361,  -14'd619,  -14'd475,  14'd678,  
-14'd104,  -14'd627,  -14'd1039,  -14'd12,  -14'd222,  -14'd1296,  -14'd630,  14'd263,  -14'd217,  14'd280,  -14'd12,  -14'd1362,  14'd340,  -14'd578,  -14'd232,  14'd797,  
-14'd875,  14'd352,  -14'd753,  14'd1320,  -14'd38,  -14'd822,  -14'd286,  -14'd326,  -14'd535,  14'd163,  14'd459,  -14'd124,  -14'd1467,  -14'd808,  -14'd356,  14'd1146,  
14'd75,  -14'd417,  -14'd713,  -14'd1178,  -14'd476,  -14'd735,  14'd175,  -14'd475,  -14'd214,  -14'd358,  -14'd78,  -14'd980,  14'd261,  14'd453,  -14'd743,  -14'd814,  
-14'd1195,  14'd327,  14'd318,  14'd888,  -14'd7,  -14'd374,  -14'd1375,  14'd186,  14'd472,  14'd797,  -14'd1523,  -14'd1685,  -14'd1089,  14'd673,  -14'd727,  -14'd542,  
-14'd1066,  -14'd351,  14'd943,  -14'd449,  14'd323,  14'd40,  14'd757,  -14'd623,  -14'd784,  -14'd530,  -14'd234,  -14'd1348,  -14'd859,  -14'd841,  14'd10,  14'd445,  
14'd143,  14'd186,  -14'd727,  -14'd952,  -14'd275,  14'd1242,  -14'd251,  -14'd423,  14'd648,  -14'd1288,  14'd107,  -14'd648,  14'd127,  -14'd413,  14'd745,  -14'd329,  
-14'd1548,  14'd84,  14'd329,  -14'd954,  -14'd480,  14'd817,  -14'd24,  14'd447,  -14'd768,  -14'd823,  -14'd1211,  14'd116,  -14'd795,  -14'd131,  -14'd786,  14'd7,  
-14'd1643,  14'd1464,  -14'd418,  -14'd866,  -14'd462,  14'd830,  14'd249,  -14'd669,  -14'd109,  -14'd248,  14'd269,  -14'd14,  -14'd965,  -14'd176,  -14'd502,  -14'd469,  
14'd633,  -14'd667,  14'd175,  -14'd298,  14'd96,  -14'd99,  -14'd193,  -14'd316,  -14'd545,  14'd112,  14'd222,  -14'd882,  -14'd1624,  -14'd89,  -14'd326,  -14'd1065,  
-14'd704,  -14'd288,  14'd45,  -14'd773,  -14'd158,  14'd384,  14'd296,  -14'd323,  14'd1266,  -14'd142,  -14'd757,  14'd1382,  14'd266,  14'd128,  -14'd895,  -14'd854,  
-14'd202,  14'd972,  14'd721,  -14'd440,  -14'd118,  14'd112,  -14'd599,  14'd600,  -14'd413,  -14'd829,  -14'd1224,  14'd796,  -14'd1521,  -14'd1754,  -14'd419,  -14'd92,  

-14'd92,  14'd426,  -14'd1259,  14'd634,  -14'd1660,  -14'd724,  -14'd1135,  -14'd883,  14'd150,  -14'd872,  14'd1284,  14'd158,  -14'd783,  -14'd1661,  -14'd813,  -14'd1211,  
-14'd250,  -14'd1417,  -14'd878,  14'd201,  -14'd21,  -14'd1194,  -14'd1298,  14'd1176,  14'd959,  14'd668,  -14'd96,  14'd494,  -14'd1210,  -14'd1498,  14'd544,  -14'd341,  
14'd373,  -14'd1369,  -14'd409,  14'd190,  -14'd360,  14'd29,  -14'd1951,  -14'd548,  -14'd1186,  14'd2107,  14'd749,  -14'd878,  14'd735,  -14'd3721,  -14'd274,  14'd42,  
-14'd1205,  -14'd3235,  -14'd1231,  14'd1568,  14'd995,  14'd917,  -14'd1238,  14'd371,  14'd1468,  14'd1274,  -14'd799,  -14'd656,  -14'd206,  -14'd1967,  -14'd1053,  14'd270,  
-14'd3067,  -14'd1677,  14'd670,  14'd337,  -14'd78,  14'd332,  14'd145,  14'd506,  -14'd772,  14'd30,  -14'd1539,  -14'd1306,  14'd627,  -14'd434,  14'd202,  -14'd2423,  
14'd382,  14'd282,  14'd31,  14'd284,  -14'd223,  14'd1586,  14'd241,  14'd145,  -14'd311,  -14'd538,  14'd1073,  14'd9,  -14'd1874,  -14'd592,  -14'd703,  14'd688,  
14'd1199,  14'd1702,  -14'd149,  14'd312,  -14'd44,  -14'd930,  14'd92,  -14'd186,  14'd1063,  14'd112,  -14'd860,  -14'd30,  14'd334,  -14'd1367,  -14'd424,  14'd969,  
14'd156,  -14'd388,  -14'd1758,  -14'd967,  -14'd341,  14'd1677,  -14'd101,  -14'd1217,  -14'd166,  -14'd400,  14'd159,  14'd1159,  14'd365,  -14'd698,  14'd349,  -14'd1,  
-14'd604,  14'd1271,  14'd687,  14'd1535,  -14'd727,  -14'd831,  14'd736,  14'd1054,  14'd2182,  14'd1858,  14'd712,  14'd576,  14'd63,  14'd150,  14'd108,  -14'd37,  
-14'd2717,  -14'd1886,  -14'd1192,  14'd251,  -14'd791,  -14'd1114,  14'd540,  14'd64,  14'd767,  -14'd1493,  14'd551,  -14'd1133,  -14'd964,  14'd141,  -14'd629,  -14'd614,  
14'd1,  14'd310,  -14'd19,  -14'd192,  14'd51,  14'd1438,  14'd928,  14'd794,  -14'd150,  14'd494,  -14'd1863,  14'd155,  14'd1072,  14'd870,  -14'd17,  -14'd132,  
-14'd460,  14'd179,  14'd685,  14'd157,  -14'd697,  -14'd699,  14'd263,  14'd477,  14'd257,  -14'd565,  -14'd348,  14'd869,  14'd352,  -14'd1264,  14'd644,  -14'd427,  
-14'd346,  14'd982,  -14'd424,  -14'd659,  14'd200,  -14'd1149,  -14'd1060,  -14'd676,  -14'd1386,  14'd241,  14'd862,  -14'd534,  14'd689,  -14'd1204,  -14'd140,  14'd600,  
14'd1823,  -14'd356,  -14'd80,  -14'd397,  14'd899,  14'd1094,  14'd487,  -14'd537,  -14'd263,  -14'd1320,  14'd1203,  14'd575,  -14'd904,  14'd653,  -14'd202,  14'd289,  
14'd822,  -14'd711,  14'd1142,  -14'd102,  14'd495,  -14'd40,  14'd956,  14'd1383,  14'd518,  -14'd1838,  14'd841,  14'd1334,  14'd126,  14'd1148,  14'd358,  14'd142,  
14'd302,  -14'd107,  14'd289,  -14'd376,  14'd1494,  14'd925,  -14'd463,  14'd18,  -14'd877,  -14'd186,  -14'd611,  14'd448,  14'd172,  14'd1580,  -14'd24,  -14'd1141,  
14'd79,  -14'd172,  -14'd1383,  -14'd71,  -14'd369,  -14'd396,  -14'd1063,  14'd1104,  14'd8,  -14'd1724,  14'd829,  -14'd1096,  14'd14,  14'd522,  14'd514,  14'd1151,  
-14'd1054,  14'd1333,  -14'd303,  -14'd1028,  14'd192,  -14'd134,  14'd162,  14'd1163,  -14'd773,  14'd56,  14'd1075,  -14'd515,  -14'd927,  14'd392,  -14'd1406,  14'd418,  
14'd1588,  14'd1579,  14'd823,  -14'd1021,  -14'd1124,  14'd346,  -14'd63,  -14'd962,  -14'd611,  14'd836,  14'd534,  14'd317,  14'd626,  14'd418,  14'd837,  -14'd695,  
14'd697,  14'd1342,  -14'd1362,  14'd75,  14'd451,  14'd381,  -14'd465,  14'd987,  -14'd1325,  -14'd877,  -14'd536,  -14'd1196,  -14'd32,  -14'd159,  14'd1037,  14'd272,  
-14'd98,  14'd1151,  -14'd189,  -14'd821,  14'd575,  -14'd513,  -14'd1292,  -14'd1462,  14'd623,  14'd625,  -14'd50,  14'd12,  -14'd1828,  -14'd380,  -14'd124,  -14'd662,  
-14'd1023,  -14'd1591,  14'd1311,  14'd326,  -14'd299,  -14'd813,  14'd459,  -14'd503,  14'd675,  14'd245,  14'd281,  -14'd144,  -14'd1476,  -14'd841,  -14'd82,  -14'd15,  
-14'd1381,  -14'd387,  14'd584,  -14'd560,  14'd172,  14'd785,  14'd1495,  -14'd1072,  14'd2062,  14'd1637,  -14'd504,  -14'd780,  -14'd1185,  14'd2152,  14'd694,  14'd244,  
-14'd763,  -14'd318,  -14'd582,  -14'd1397,  14'd158,  14'd1093,  -14'd1203,  14'd166,  14'd562,  14'd478,  14'd148,  14'd6,  14'd533,  14'd794,  14'd235,  -14'd1128,  
-14'd1054,  -14'd997,  14'd369,  14'd1278,  -14'd1623,  -14'd191,  -14'd816,  14'd43,  14'd132,  14'd338,  -14'd1015,  -14'd506,  14'd105,  -14'd1795,  14'd801,  -14'd1112,  

-14'd243,  -14'd69,  -14'd1079,  14'd420,  14'd327,  -14'd567,  -14'd221,  14'd416,  -14'd1220,  -14'd955,  -14'd1235,  14'd470,  -14'd466,  14'd132,  14'd473,  -14'd2056,  
14'd168,  14'd1443,  -14'd1116,  -14'd512,  14'd1416,  -14'd25,  -14'd1290,  -14'd552,  14'd418,  14'd532,  -14'd638,  14'd532,  -14'd400,  -14'd983,  14'd247,  -14'd361,  
-14'd376,  14'd1254,  -14'd1505,  -14'd396,  14'd636,  14'd439,  14'd1523,  -14'd566,  -14'd1165,  14'd595,  14'd524,  14'd874,  -14'd182,  -14'd1121,  -14'd506,  14'd595,  
-14'd1396,  -14'd378,  14'd574,  -14'd1202,  14'd1288,  -14'd1238,  14'd138,  -14'd1379,  14'd732,  -14'd831,  -14'd1388,  14'd1318,  14'd286,  14'd720,  -14'd765,  14'd1098,  
-14'd1197,  -14'd1927,  -14'd690,  -14'd1198,  -14'd820,  -14'd180,  -14'd731,  -14'd258,  -14'd97,  -14'd892,  -14'd350,  -14'd1419,  -14'd569,  14'd267,  -14'd1008,  -14'd466,  
14'd252,  14'd322,  -14'd171,  14'd834,  -14'd212,  14'd217,  14'd71,  -14'd206,  14'd1648,  -14'd484,  -14'd119,  14'd218,  14'd452,  14'd853,  -14'd1047,  -14'd780,  
14'd880,  14'd7,  -14'd306,  -14'd1015,  -14'd1251,  14'd271,  -14'd442,  14'd790,  -14'd1014,  -14'd457,  -14'd728,  -14'd543,  14'd959,  -14'd478,  -14'd853,  14'd1055,  
14'd1559,  -14'd1,  -14'd191,  -14'd264,  -14'd946,  -14'd534,  14'd509,  14'd1548,  -14'd755,  -14'd531,  -14'd839,  14'd1125,  14'd905,  14'd517,  14'd1639,  14'd247,  
-14'd33,  -14'd187,  14'd113,  -14'd260,  14'd42,  14'd351,  14'd2134,  -14'd818,  14'd411,  -14'd522,  -14'd51,  14'd1925,  14'd388,  14'd2818,  14'd238,  -14'd428,  
-14'd1153,  14'd42,  -14'd543,  -14'd446,  14'd233,  14'd260,  14'd879,  14'd944,  -14'd399,  14'd593,  -14'd128,  -14'd1618,  -14'd228,  14'd663,  -14'd607,  -14'd1775,  
-14'd179,  -14'd8,  -14'd339,  -14'd197,  14'd1434,  14'd306,  -14'd253,  -14'd491,  -14'd239,  14'd296,  -14'd1803,  -14'd458,  -14'd1233,  14'd1142,  -14'd1133,  -14'd535,  
14'd616,  14'd228,  14'd1811,  14'd884,  14'd1243,  -14'd88,  -14'd1097,  -14'd659,  -14'd402,  -14'd1401,  14'd233,  14'd1140,  14'd159,  -14'd861,  14'd429,  -14'd457,  
14'd468,  14'd555,  14'd397,  -14'd1029,  -14'd1412,  14'd1639,  -14'd833,  14'd1412,  14'd476,  -14'd938,  14'd1875,  14'd434,  14'd543,  14'd395,  -14'd1155,  14'd1419,  
-14'd1107,  -14'd5,  14'd888,  14'd1186,  -14'd1396,  -14'd677,  14'd728,  14'd378,  14'd787,  -14'd468,  14'd731,  -14'd585,  14'd476,  14'd781,  14'd727,  -14'd572,  
14'd506,  -14'd892,  -14'd86,  14'd32,  14'd145,  -14'd1057,  -14'd793,  -14'd429,  14'd520,  -14'd1197,  -14'd76,  -14'd1955,  14'd898,  14'd981,  -14'd525,  -14'd1424,  
-14'd823,  -14'd408,  -14'd1409,  14'd276,  -14'd1282,  14'd776,  -14'd338,  -14'd726,  -14'd253,  14'd644,  -14'd332,  -14'd1347,  -14'd245,  14'd78,  -14'd1049,  14'd549,  
-14'd177,  14'd109,  -14'd783,  14'd900,  -14'd275,  -14'd135,  -14'd743,  14'd1453,  14'd619,  -14'd1350,  14'd1773,  -14'd872,  14'd142,  14'd23,  14'd198,  14'd61,  
14'd551,  -14'd388,  14'd1587,  -14'd417,  14'd1193,  -14'd1151,  -14'd468,  -14'd234,  14'd1335,  14'd1432,  14'd637,  14'd433,  14'd793,  -14'd64,  -14'd1626,  -14'd534,  
14'd932,  -14'd499,  14'd230,  -14'd328,  -14'd1026,  14'd486,  -14'd31,  14'd454,  14'd936,  14'd31,  14'd259,  -14'd425,  -14'd374,  14'd1274,  14'd129,  -14'd1374,  
14'd611,  -14'd1401,  -14'd2193,  -14'd1241,  -14'd1195,  -14'd1148,  -14'd295,  -14'd1182,  -14'd1864,  14'd1351,  -14'd783,  -14'd353,  14'd172,  14'd453,  -14'd125,  -14'd1582,  
14'd215,  14'd60,  14'd118,  -14'd436,  14'd1139,  -14'd374,  14'd1199,  -14'd1405,  -14'd1553,  14'd799,  14'd1371,  14'd476,  -14'd858,  14'd669,  -14'd38,  14'd1216,  
-14'd169,  14'd207,  -14'd811,  14'd433,  14'd179,  -14'd692,  14'd1461,  -14'd28,  14'd2166,  -14'd1,  14'd676,  -14'd893,  -14'd1508,  -14'd263,  14'd165,  14'd950,  
-14'd257,  14'd203,  14'd766,  -14'd455,  14'd871,  -14'd603,  -14'd1384,  -14'd247,  14'd209,  -14'd1083,  -14'd1856,  -14'd269,  14'd257,  14'd2131,  14'd236,  14'd258,  
-14'd388,  14'd150,  -14'd149,  14'd415,  -14'd557,  14'd679,  -14'd1071,  -14'd913,  -14'd323,  14'd1135,  -14'd118,  -14'd130,  -14'd1504,  -14'd43,  14'd1578,  14'd1317,  
-14'd1918,  14'd417,  14'd1363,  14'd160,  14'd138,  14'd1453,  14'd1127,  -14'd1425,  14'd92,  14'd2931,  14'd996,  -14'd1287,  -14'd294,  -14'd1168,  14'd756,  -14'd592,  

-14'd1485,  14'd823,  -14'd403,  14'd1263,  -14'd206,  14'd431,  -14'd183,  -14'd967,  14'd944,  -14'd21,  14'd212,  14'd946,  14'd400,  14'd306,  14'd80,  14'd115,  
-14'd763,  14'd1230,  14'd195,  14'd1374,  -14'd145,  -14'd193,  -14'd812,  14'd1657,  -14'd1327,  14'd209,  -14'd821,  14'd1365,  -14'd299,  14'd1002,  -14'd380,  14'd918,  
-14'd758,  -14'd1795,  14'd1484,  -14'd1040,  14'd329,  14'd214,  14'd613,  -14'd465,  14'd1750,  14'd91,  -14'd361,  -14'd1129,  14'd763,  14'd2372,  14'd532,  -14'd350,  
-14'd769,  -14'd1818,  -14'd1099,  14'd33,  -14'd913,  14'd354,  14'd318,  -14'd64,  -14'd910,  -14'd136,  14'd992,  14'd1306,  -14'd816,  -14'd1087,  -14'd468,  -14'd554,  
-14'd529,  -14'd1149,  -14'd960,  -14'd282,  -14'd736,  -14'd169,  14'd1532,  -14'd138,  -14'd1370,  -14'd1552,  14'd109,  -14'd539,  -14'd381,  14'd659,  14'd42,  14'd436,  
-14'd793,  14'd515,  -14'd550,  -14'd633,  -14'd660,  14'd82,  -14'd741,  14'd67,  -14'd1575,  -14'd615,  14'd713,  14'd94,  14'd585,  14'd1371,  -14'd258,  14'd122,  
14'd936,  -14'd1085,  14'd526,  14'd65,  -14'd173,  -14'd464,  14'd433,  -14'd702,  -14'd1250,  -14'd47,  -14'd38,  14'd183,  -14'd1076,  -14'd100,  14'd383,  14'd800,  
14'd46,  -14'd1377,  -14'd279,  14'd58,  -14'd530,  -14'd526,  -14'd270,  14'd1020,  14'd1274,  -14'd985,  14'd281,  -14'd226,  -14'd17,  -14'd223,  14'd1047,  14'd845,  
-14'd377,  -14'd1828,  14'd5,  14'd250,  -14'd971,  -14'd320,  -14'd137,  14'd537,  -14'd218,  -14'd206,  14'd44,  -14'd347,  -14'd147,  -14'd216,  14'd376,  -14'd1269,  
-14'd1169,  14'd332,  -14'd1480,  -14'd240,  -14'd1827,  14'd1613,  -14'd863,  14'd392,  14'd522,  -14'd650,  14'd638,  -14'd614,  14'd481,  -14'd124,  -14'd301,  14'd1424,  
-14'd567,  -14'd493,  14'd237,  14'd203,  -14'd1403,  -14'd1579,  -14'd1838,  14'd61,  14'd640,  14'd1421,  14'd117,  -14'd548,  -14'd89,  -14'd235,  -14'd103,  -14'd202,  
14'd843,  -14'd1213,  14'd995,  14'd62,  -14'd2010,  14'd151,  -14'd2909,  14'd414,  -14'd2012,  14'd2174,  -14'd225,  14'd751,  -14'd466,  -14'd395,  14'd681,  14'd1415,  
-14'd815,  -14'd851,  -14'd686,  -14'd419,  14'd831,  -14'd665,  -14'd1526,  -14'd411,  -14'd2082,  -14'd367,  -14'd390,  -14'd273,  14'd443,  14'd527,  14'd1079,  14'd821,  
-14'd260,  14'd622,  -14'd1247,  -14'd146,  14'd452,  -14'd1368,  -14'd629,  14'd430,  -14'd756,  -14'd1234,  14'd74,  14'd870,  -14'd1000,  -14'd1065,  -14'd665,  -14'd76,  
-14'd3689,  -14'd1864,  14'd165,  -14'd628,  14'd1073,  -14'd765,  -14'd1281,  -14'd312,  14'd22,  14'd1634,  -14'd732,  14'd651,  -14'd1560,  -14'd625,  -14'd179,  -14'd1765,  
-14'd2299,  -14'd2012,  -14'd349,  14'd1722,  -14'd296,  -14'd415,  -14'd3541,  14'd867,  14'd814,  14'd332,  14'd180,  -14'd767,  14'd157,  -14'd742,  -14'd232,  -14'd1097,  
-14'd1702,  -14'd1323,  14'd1942,  -14'd948,  14'd738,  -14'd510,  -14'd1504,  -14'd823,  -14'd707,  14'd1447,  14'd952,  14'd355,  -14'd205,  -14'd558,  -14'd1080,  -14'd316,  
14'd652,  -14'd1198,  14'd562,  14'd179,  -14'd725,  14'd647,  14'd763,  14'd522,  14'd660,  14'd329,  14'd588,  14'd471,  -14'd246,  -14'd497,  14'd80,  -14'd251,  
-14'd461,  -14'd3,  -14'd733,  14'd1461,  14'd628,  14'd1408,  14'd336,  14'd1256,  -14'd87,  -14'd931,  14'd1084,  14'd1107,  14'd742,  14'd919,  14'd1736,  14'd1562,  
-14'd501,  -14'd386,  -14'd58,  14'd909,  -14'd141,  14'd327,  14'd1200,  14'd1060,  14'd1842,  14'd1053,  -14'd230,  14'd106,  -14'd1060,  14'd636,  14'd820,  14'd282,  
-14'd1036,  14'd205,  -14'd1509,  14'd1030,  14'd175,  14'd1102,  -14'd74,  14'd571,  14'd3588,  14'd1131,  14'd1235,  14'd1628,  -14'd404,  -14'd1050,  14'd760,  14'd336,  
-14'd298,  -14'd107,  -14'd471,  14'd1624,  14'd787,  14'd186,  14'd5,  14'd511,  14'd893,  14'd364,  14'd469,  14'd678,  14'd1511,  -14'd4308,  14'd392,  14'd1111,  
14'd1123,  14'd882,  -14'd1131,  -14'd538,  14'd821,  14'd498,  -14'd623,  14'd893,  14'd966,  14'd752,  14'd285,  14'd122,  14'd2051,  -14'd1337,  -14'd126,  -14'd76,  
14'd1762,  14'd980,  -14'd505,  -14'd488,  14'd86,  14'd629,  14'd708,  14'd1093,  14'd862,  -14'd148,  -14'd510,  -14'd822,  14'd1162,  14'd254,  -14'd313,  14'd480,  
14'd1460,  14'd2064,  14'd44,  14'd728,  -14'd964,  14'd937,  -14'd682,  14'd115,  14'd845,  -14'd622,  -14'd673,  14'd217,  14'd989,  14'd928,  14'd511,  14'd335,  

-14'd520,  14'd237,  14'd500,  14'd790,  -14'd786,  -14'd130,  -14'd182,  14'd19,  -14'd466,  14'd955,  14'd874,  -14'd760,  14'd872,  -14'd261,  -14'd133,  14'd927,  
14'd252,  14'd212,  14'd828,  -14'd669,  -14'd167,  -14'd304,  -14'd1677,  -14'd991,  14'd1497,  -14'd111,  -14'd621,  -14'd664,  14'd427,  -14'd860,  14'd118,  -14'd397,  
-14'd242,  14'd369,  14'd811,  -14'd886,  -14'd134,  14'd500,  -14'd751,  14'd129,  14'd177,  14'd1027,  14'd442,  -14'd477,  -14'd1255,  14'd317,  -14'd3,  -14'd1538,  
-14'd865,  -14'd958,  -14'd608,  14'd80,  14'd803,  -14'd242,  14'd192,  -14'd546,  14'd157,  -14'd32,  -14'd132,  14'd1012,  14'd10,  -14'd683,  14'd257,  -14'd1554,  
14'd630,  14'd320,  -14'd853,  -14'd185,  -14'd324,  14'd190,  -14'd1634,  -14'd853,  14'd620,  -14'd748,  14'd1025,  -14'd103,  14'd641,  -14'd163,  14'd599,  -14'd189,  
-14'd722,  14'd873,  14'd243,  14'd41,  14'd133,  -14'd1288,  -14'd1048,  14'd153,  -14'd498,  14'd498,  14'd1167,  -14'd626,  14'd1283,  14'd129,  -14'd664,  14'd763,  
14'd1399,  -14'd1220,  -14'd705,  -14'd637,  -14'd682,  -14'd339,  14'd460,  14'd990,  -14'd595,  -14'd101,  -14'd1405,  -14'd1116,  -14'd510,  14'd652,  -14'd303,  -14'd322,  
14'd583,  -14'd531,  -14'd214,  -14'd943,  -14'd1192,  -14'd414,  14'd299,  14'd436,  -14'd1614,  14'd115,  -14'd1248,  -14'd1262,  14'd257,  -14'd766,  -14'd1024,  -14'd1126,  
-14'd277,  14'd314,  -14'd787,  14'd57,  -14'd1835,  14'd319,  14'd369,  -14'd177,  -14'd436,  -14'd860,  14'd842,  -14'd1048,  14'd92,  -14'd89,  14'd395,  14'd207,  
-14'd423,  14'd1083,  -14'd999,  14'd522,  -14'd948,  -14'd443,  -14'd846,  -14'd614,  -14'd1602,  -14'd34,  14'd1318,  14'd627,  14'd173,  14'd78,  -14'd1634,  14'd393,  
14'd389,  -14'd585,  -14'd1575,  -14'd1381,  14'd82,  -14'd180,  -14'd785,  -14'd989,  14'd57,  14'd487,  -14'd344,  14'd23,  -14'd1361,  -14'd1363,  14'd98,  14'd785,  
-14'd1435,  -14'd1205,  14'd1020,  14'd92,  -14'd433,  -14'd1178,  14'd1185,  -14'd604,  14'd597,  -14'd210,  14'd1040,  14'd233,  14'd658,  14'd103,  -14'd1109,  -14'd1284,  
-14'd410,  14'd335,  14'd144,  -14'd87,  14'd601,  14'd1034,  -14'd917,  -14'd563,  -14'd930,  14'd1153,  14'd172,  14'd282,  14'd155,  -14'd248,  -14'd645,  -14'd415,  
-14'd612,  -14'd242,  14'd282,  -14'd962,  -14'd635,  14'd978,  -14'd1517,  14'd851,  -14'd1350,  -14'd266,  14'd222,  14'd346,  14'd465,  -14'd275,  -14'd496,  -14'd57,  
-14'd265,  -14'd1320,  -14'd339,  14'd180,  14'd734,  14'd804,  -14'd1390,  -14'd765,  14'd600,  14'd959,  -14'd520,  -14'd79,  -14'd1187,  14'd283,  14'd646,  -14'd734,  
-14'd621,  -14'd23,  14'd702,  14'd659,  14'd585,  14'd912,  14'd276,  -14'd1243,  -14'd724,  -14'd606,  -14'd1246,  -14'd564,  14'd416,  -14'd1023,  -14'd968,  14'd1274,  
14'd782,  14'd1279,  14'd429,  -14'd145,  -14'd761,  -14'd362,  -14'd425,  -14'd496,  -14'd1163,  -14'd648,  -14'd173,  -14'd1123,  -14'd512,  14'd277,  14'd1228,  14'd384,  
-14'd668,  14'd463,  -14'd93,  -14'd1053,  -14'd1189,  14'd702,  14'd179,  -14'd143,  14'd434,  -14'd316,  14'd58,  14'd410,  -14'd522,  14'd461,  -14'd267,  -14'd4,  
14'd526,  -14'd580,  -14'd939,  14'd412,  14'd51,  -14'd52,  -14'd353,  14'd424,  14'd1399,  -14'd170,  14'd516,  -14'd656,  -14'd103,  14'd533,  -14'd31,  -14'd583,  
-14'd201,  -14'd1252,  -14'd293,  -14'd381,  14'd459,  14'd449,  -14'd627,  14'd473,  -14'd200,  14'd594,  -14'd706,  14'd683,  14'd305,  -14'd716,  14'd416,  -14'd810,  
14'd29,  14'd528,  14'd1559,  -14'd1509,  14'd302,  -14'd531,  14'd1119,  14'd90,  14'd998,  14'd486,  -14'd483,  14'd354,  14'd1490,  -14'd797,  -14'd198,  -14'd300,  
-14'd823,  -14'd65,  -14'd145,  14'd513,  14'd737,  -14'd1438,  14'd689,  -14'd1081,  -14'd1186,  14'd952,  -14'd816,  -14'd48,  14'd526,  -14'd87,  14'd99,  -14'd130,  
-14'd1154,  14'd302,  -14'd239,  -14'd1234,  14'd745,  -14'd1231,  14'd67,  14'd1020,  -14'd596,  -14'd67,  -14'd262,  14'd803,  14'd440,  -14'd28,  -14'd716,  14'd52,  
14'd335,  14'd229,  -14'd1000,  14'd1076,  14'd610,  -14'd612,  -14'd1429,  -14'd185,  14'd1225,  14'd1169,  -14'd634,  14'd486,  -14'd886,  -14'd592,  14'd844,  14'd940,  
-14'd1341,  14'd337,  -14'd309,  14'd664,  -14'd50,  14'd309,  14'd882,  14'd1363,  -14'd47,  -14'd798,  14'd842,  14'd618,  14'd478,  14'd251,  -14'd429,  14'd708,  

14'd27,  14'd72,  -14'd1623,  14'd329,  14'd677,  -14'd116,  14'd1030,  14'd1118,  14'd394,  -14'd1304,  14'd1622,  14'd573,  14'd2015,  14'd395,  14'd1039,  14'd1772,  
14'd74,  14'd1199,  -14'd1758,  14'd904,  14'd261,  14'd935,  14'd308,  14'd882,  14'd1092,  14'd380,  14'd1401,  -14'd412,  14'd843,  -14'd1809,  14'd1255,  14'd577,  
-14'd2124,  -14'd436,  14'd434,  -14'd609,  14'd951,  14'd537,  -14'd2588,  -14'd75,  -14'd1358,  -14'd1788,  -14'd1476,  -14'd408,  14'd1485,  14'd936,  14'd270,  14'd1297,  
-14'd39,  -14'd1371,  -14'd834,  -14'd1004,  -14'd1048,  -14'd656,  14'd319,  14'd353,  -14'd555,  14'd740,  14'd525,  14'd569,  -14'd1481,  -14'd716,  -14'd771,  -14'd2564,  
-14'd8,  -14'd1085,  -14'd209,  -14'd1515,  -14'd1697,  14'd160,  -14'd419,  -14'd84,  -14'd20,  -14'd223,  -14'd892,  -14'd34,  -14'd1500,  14'd1317,  -14'd2031,  -14'd859,  
-14'd1118,  14'd1093,  14'd194,  -14'd249,  14'd570,  14'd651,  14'd1920,  -14'd470,  14'd183,  -14'd147,  14'd1468,  14'd253,  -14'd1233,  -14'd528,  -14'd1453,  -14'd986,  
14'd233,  -14'd141,  -14'd142,  14'd3,  14'd824,  14'd530,  14'd7,  14'd9,  14'd857,  14'd1123,  14'd821,  -14'd564,  -14'd114,  -14'd525,  14'd1070,  -14'd861,  
14'd80,  14'd91,  14'd144,  -14'd298,  14'd1058,  -14'd835,  -14'd1258,  14'd296,  -14'd1126,  -14'd110,  -14'd104,  14'd441,  -14'd717,  14'd830,  14'd14,  14'd320,  
-14'd88,  -14'd1271,  -14'd1728,  -14'd718,  -14'd530,  -14'd1796,  -14'd624,  -14'd1610,  14'd1012,  -14'd1130,  -14'd1235,  -14'd990,  -14'd2184,  14'd1004,  -14'd670,  -14'd695,  
-14'd1899,  14'd479,  14'd743,  -14'd707,  -14'd779,  -14'd461,  -14'd774,  -14'd2049,  -14'd1970,  14'd677,  -14'd954,  14'd223,  -14'd2257,  14'd2128,  -14'd807,  -14'd433,  
-14'd340,  -14'd189,  -14'd1463,  -14'd294,  14'd295,  14'd89,  14'd1462,  -14'd1540,  14'd228,  -14'd944,  -14'd648,  -14'd1494,  -14'd4,  14'd143,  -14'd818,  14'd236,  
-14'd571,  14'd975,  -14'd366,  -14'd81,  14'd386,  -14'd0,  -14'd431,  14'd28,  14'd2143,  14'd743,  -14'd911,  -14'd158,  14'd592,  -14'd317,  14'd1074,  14'd1075,  
-14'd90,  14'd658,  14'd49,  -14'd36,  -14'd526,  14'd580,  -14'd256,  -14'd120,  14'd1775,  14'd903,  14'd997,  -14'd555,  14'd693,  14'd769,  -14'd791,  -14'd258,  
-14'd2308,  14'd846,  -14'd2426,  14'd2121,  14'd38,  14'd889,  14'd856,  -14'd306,  14'd1987,  -14'd1185,  14'd2923,  14'd478,  -14'd302,  14'd275,  -14'd691,  14'd961,  
-14'd2099,  -14'd149,  14'd1646,  14'd1649,  -14'd252,  -14'd303,  -14'd124,  14'd597,  -14'd405,  -14'd268,  14'd3263,  14'd158,  14'd1918,  -14'd486,  14'd55,  14'd881,  
14'd2221,  14'd435,  14'd1144,  -14'd973,  -14'd1406,  14'd1233,  -14'd788,  -14'd230,  14'd127,  14'd147,  -14'd2147,  -14'd1038,  -14'd1396,  14'd1682,  14'd481,  -14'd1882,  
14'd800,  -14'd200,  -14'd54,  -14'd384,  -14'd87,  -14'd1476,  -14'd890,  -14'd576,  -14'd456,  -14'd146,  -14'd724,  -14'd392,  14'd375,  14'd935,  14'd2077,  14'd1341,  
14'd606,  -14'd1212,  14'd439,  -14'd1501,  14'd996,  14'd87,  14'd978,  -14'd1377,  14'd259,  14'd1400,  14'd1347,  14'd144,  -14'd355,  -14'd380,  -14'd606,  14'd396,  
-14'd24,  14'd2955,  -14'd926,  14'd688,  14'd451,  -14'd306,  14'd76,  14'd184,  14'd677,  -14'd1194,  14'd1598,  -14'd174,  14'd750,  14'd226,  14'd811,  14'd1176,  
-14'd220,  -14'd821,  -14'd842,  14'd44,  14'd71,  -14'd1494,  -14'd76,  -14'd917,  -14'd1353,  14'd971,  14'd1629,  -14'd1331,  -14'd81,  14'd97,  14'd268,  14'd2207,  
14'd348,  14'd646,  14'd1533,  14'd1409,  -14'd1022,  14'd658,  -14'd1609,  14'd951,  -14'd1860,  -14'd176,  -14'd1634,  -14'd1339,  -14'd1052,  14'd1249,  14'd280,  -14'd1955,  
14'd893,  -14'd540,  -14'd847,  -14'd469,  -14'd846,  14'd29,  -14'd112,  -14'd214,  -14'd1262,  -14'd546,  14'd18,  -14'd1334,  14'd423,  14'd1271,  14'd851,  14'd191,  
14'd521,  -14'd355,  -14'd323,  14'd648,  14'd2086,  -14'd808,  14'd1477,  14'd1262,  -14'd1411,  -14'd1757,  -14'd267,  -14'd1325,  -14'd954,  -14'd735,  -14'd1304,  14'd96,  
-14'd2318,  14'd1279,  14'd240,  -14'd266,  14'd115,  14'd542,  -14'd907,  14'd1372,  -14'd242,  14'd935,  -14'd1194,  -14'd1992,  -14'd1171,  14'd1229,  -14'd1793,  14'd53,  
-14'd2307,  -14'd373,  14'd116,  14'd1681,  14'd599,  -14'd266,  -14'd686,  -14'd231,  -14'd1695,  14'd2808,  14'd211,  -14'd488,  -14'd410,  -14'd232,  -14'd119,  14'd455,  

-14'd1218,  -14'd457,  -14'd540,  -14'd258,  14'd1098,  -14'd385,  14'd507,  14'd944,  -14'd358,  14'd27,  14'd1333,  -14'd1677,  -14'd56,  -14'd1410,  14'd1251,  14'd193,  
-14'd1243,  -14'd369,  -14'd11,  14'd403,  14'd531,  -14'd305,  -14'd2760,  -14'd45,  -14'd1503,  14'd1338,  -14'd1964,  -14'd738,  14'd994,  -14'd2508,  -14'd42,  14'd28,  
-14'd388,  -14'd1514,  14'd1115,  14'd1795,  -14'd889,  14'd431,  14'd1160,  14'd1371,  -14'd639,  14'd1261,  14'd1242,  -14'd612,  -14'd1109,  -14'd1872,  14'd413,  14'd1422,  
14'd1576,  -14'd2470,  -14'd935,  14'd771,  -14'd86,  14'd1591,  14'd1417,  14'd882,  14'd1020,  -14'd606,  14'd293,  14'd765,  14'd1244,  14'd2165,  -14'd555,  -14'd770,  
-14'd1713,  -14'd57,  14'd566,  -14'd1037,  14'd535,  14'd850,  14'd272,  -14'd749,  14'd1609,  -14'd1092,  14'd642,  14'd647,  -14'd2148,  14'd859,  -14'd182,  -14'd520,  
-14'd1697,  14'd100,  -14'd1364,  -14'd636,  -14'd835,  -14'd1681,  -14'd2010,  -14'd88,  -14'd507,  -14'd1286,  14'd1433,  -14'd64,  -14'd520,  -14'd852,  -14'd24,  14'd657,  
-14'd693,  -14'd1041,  -14'd1704,  -14'd1571,  14'd1083,  14'd236,  -14'd386,  14'd392,  -14'd393,  -14'd187,  14'd1257,  14'd100,  -14'd676,  -14'd1116,  14'd587,  14'd525,  
14'd898,  -14'd568,  -14'd1114,  14'd562,  -14'd5,  -14'd448,  -14'd102,  -14'd80,  -14'd1324,  14'd1073,  -14'd118,  -14'd13,  -14'd411,  -14'd1714,  14'd1178,  14'd1095,  
14'd2081,  14'd195,  -14'd635,  -14'd163,  -14'd284,  -14'd928,  14'd1436,  14'd911,  -14'd447,  14'd529,  -14'd401,  14'd154,  -14'd720,  14'd249,  14'd270,  14'd325,  
-14'd601,  14'd935,  -14'd328,  14'd1091,  -14'd874,  14'd1064,  14'd541,  -14'd398,  -14'd1494,  -14'd42,  14'd189,  -14'd963,  14'd428,  14'd347,  -14'd674,  -14'd926,  
-14'd1306,  -14'd434,  14'd249,  -14'd535,  -14'd1471,  -14'd957,  14'd1193,  14'd846,  14'd1355,  -14'd766,  14'd1042,  -14'd556,  -14'd1228,  -14'd383,  14'd317,  -14'd1306,  
14'd1034,  -14'd962,  14'd470,  -14'd945,  -14'd1874,  -14'd1500,  14'd459,  -14'd413,  -14'd280,  14'd723,  -14'd1354,  -14'd1103,  14'd250,  14'd1164,  14'd1577,  -14'd1083,  
14'd889,  -14'd453,  14'd1195,  -14'd775,  -14'd1293,  14'd302,  14'd223,  14'd305,  14'd281,  14'd269,  14'd88,  14'd748,  -14'd412,  14'd247,  -14'd624,  -14'd550,  
-14'd680,  -14'd144,  -14'd216,  14'd676,  14'd349,  14'd583,  14'd414,  14'd940,  14'd517,  14'd886,  14'd172,  14'd1136,  -14'd319,  -14'd615,  14'd74,  14'd896,  
-14'd594,  -14'd58,  14'd368,  14'd314,  -14'd383,  -14'd507,  14'd484,  -14'd200,  14'd275,  14'd1191,  14'd373,  -14'd782,  -14'd71,  -14'd257,  -14'd209,  -14'd868,  
-14'd1384,  -14'd1348,  14'd816,  14'd1703,  -14'd88,  14'd1215,  -14'd866,  14'd982,  14'd771,  14'd362,  14'd797,  -14'd361,  -14'd759,  14'd149,  14'd266,  14'd446,  
-14'd1980,  -14'd559,  -14'd386,  14'd337,  14'd5,  -14'd851,  14'd919,  -14'd1295,  -14'd823,  14'd1727,  14'd1253,  -14'd638,  -14'd854,  -14'd141,  14'd1283,  -14'd430,  
-14'd211,  14'd844,  14'd429,  14'd542,  -14'd119,  14'd578,  14'd305,  14'd530,  -14'd488,  -14'd1007,  -14'd1055,  -14'd102,  -14'd26,  14'd356,  -14'd244,  -14'd1080,  
14'd5,  -14'd184,  14'd1254,  14'd1464,  -14'd1686,  -14'd567,  -14'd33,  -14'd648,  -14'd1555,  -14'd981,  -14'd323,  14'd352,  14'd537,  -14'd58,  14'd150,  14'd1293,  
14'd38,  14'd337,  14'd297,  14'd426,  -14'd745,  -14'd387,  14'd867,  14'd105,  -14'd938,  -14'd235,  14'd1252,  -14'd644,  -14'd1085,  14'd659,  -14'd1350,  14'd707,  
-14'd810,  14'd703,  -14'd667,  14'd1275,  -14'd589,  -14'd210,  14'd612,  14'd105,  14'd1016,  14'd315,  14'd845,  -14'd489,  14'd644,  -14'd1687,  -14'd392,  -14'd245,  
14'd315,  14'd1058,  14'd661,  -14'd358,  14'd54,  14'd562,  -14'd382,  -14'd1501,  14'd829,  14'd842,  14'd358,  14'd1093,  14'd366,  -14'd1284,  -14'd76,  14'd315,  
14'd58,  14'd475,  14'd444,  14'd897,  -14'd521,  14'd228,  14'd87,  -14'd252,  14'd1799,  14'd124,  14'd507,  -14'd1339,  14'd885,  -14'd39,  14'd1189,  14'd179,  
14'd1508,  -14'd304,  -14'd525,  -14'd9,  -14'd451,  14'd201,  14'd1192,  -14'd63,  -14'd582,  -14'd386,  14'd1555,  -14'd597,  14'd895,  14'd1076,  -14'd1305,  -14'd1018,  
14'd540,  14'd564,  -14'd1073,  -14'd67,  14'd253,  -14'd139,  -14'd519,  -14'd36,  14'd629,  -14'd526,  14'd521,  -14'd92,  -14'd982,  -14'd84,  -14'd294,  -14'd708,  

-14'd522,  14'd1738,  14'd1372,  14'd417,  -14'd408,  14'd621,  14'd630,  -14'd1784,  14'd811,  -14'd1189,  -14'd1762,  14'd763,  -14'd772,  14'd770,  -14'd687,  -14'd550,  
-14'd183,  -14'd108,  14'd2144,  -14'd1944,  14'd230,  -14'd439,  -14'd196,  -14'd37,  14'd373,  -14'd363,  14'd380,  -14'd755,  14'd121,  14'd2335,  14'd91,  -14'd941,  
-14'd1892,  14'd433,  14'd703,  -14'd139,  -14'd728,  14'd396,  -14'd478,  14'd71,  14'd146,  -14'd929,  14'd689,  14'd481,  -14'd1658,  14'd2344,  -14'd306,  -14'd1561,  
14'd356,  14'd20,  -14'd1007,  14'd576,  -14'd261,  14'd1198,  14'd480,  -14'd327,  14'd526,  14'd738,  -14'd1410,  14'd478,  -14'd947,  14'd755,  -14'd1000,  -14'd119,  
14'd1148,  14'd589,  -14'd238,  14'd877,  -14'd486,  14'd245,  14'd978,  14'd48,  14'd1346,  -14'd685,  -14'd156,  14'd724,  14'd1170,  14'd1137,  14'd84,  14'd1041,  
14'd178,  14'd1384,  14'd184,  14'd317,  -14'd1245,  -14'd611,  14'd861,  14'd1084,  -14'd766,  14'd1867,  -14'd597,  14'd569,  -14'd689,  14'd1864,  14'd1123,  14'd482,  
14'd671,  14'd102,  14'd1814,  -14'd1127,  -14'd613,  -14'd1591,  -14'd1195,  14'd528,  14'd1147,  -14'd158,  -14'd275,  -14'd774,  14'd1069,  14'd2122,  14'd1103,  14'd1185,  
14'd139,  -14'd1244,  14'd1310,  -14'd49,  -14'd55,  -14'd91,  -14'd1113,  14'd577,  14'd1039,  14'd197,  14'd701,  -14'd676,  -14'd449,  14'd154,  -14'd1341,  -14'd1270,  
-14'd804,  14'd695,  14'd1063,  -14'd480,  14'd250,  14'd1139,  -14'd544,  14'd203,  -14'd128,  14'd825,  -14'd924,  14'd829,  -14'd662,  -14'd366,  14'd288,  14'd431,  
14'd1161,  -14'd1102,  -14'd807,  14'd96,  -14'd380,  14'd664,  -14'd323,  -14'd1259,  14'd598,  -14'd2031,  -14'd511,  -14'd464,  -14'd1285,  14'd386,  -14'd554,  14'd728,  
14'd1628,  -14'd260,  -14'd38,  14'd1656,  -14'd702,  14'd2489,  -14'd1623,  14'd745,  14'd617,  14'd153,  14'd1040,  -14'd458,  14'd2396,  14'd799,  -14'd251,  14'd694,  
-14'd441,  14'd1417,  14'd240,  14'd694,  -14'd1083,  14'd1341,  -14'd289,  14'd1731,  14'd591,  14'd1124,  -14'd199,  -14'd246,  14'd510,  -14'd699,  14'd202,  -14'd1456,  
14'd614,  -14'd161,  -14'd58,  14'd1084,  -14'd283,  14'd1626,  14'd601,  14'd555,  -14'd134,  -14'd419,  14'd1700,  14'd62,  14'd1559,  -14'd1676,  -14'd843,  14'd45,  
-14'd112,  14'd272,  -14'd950,  14'd192,  14'd81,  -14'd935,  -14'd519,  -14'd923,  -14'd15,  -14'd1162,  14'd1585,  14'd841,  14'd63,  -14'd270,  14'd268,  -14'd313,  
-14'd495,  -14'd1080,  -14'd180,  -14'd386,  -14'd439,  14'd99,  14'd725,  14'd629,  -14'd793,  -14'd942,  -14'd822,  -14'd74,  14'd2175,  -14'd259,  -14'd257,  14'd1837,  
14'd466,  14'd1582,  -14'd674,  14'd38,  14'd2971,  14'd603,  -14'd539,  -14'd758,  -14'd585,  14'd555,  -14'd234,  14'd1707,  14'd824,  -14'd224,  14'd311,  14'd1575,  
-14'd1461,  -14'd214,  -14'd291,  -14'd48,  14'd702,  -14'd1915,  14'd570,  14'd506,  -14'd299,  14'd321,  14'd330,  14'd325,  14'd422,  -14'd1144,  -14'd575,  14'd404,  
-14'd226,  -14'd1022,  14'd720,  14'd515,  14'd976,  -14'd582,  14'd576,  -14'd1326,  14'd804,  14'd107,  -14'd417,  14'd320,  -14'd172,  14'd412,  -14'd1107,  14'd107,  
14'd1320,  14'd392,  14'd862,  14'd726,  -14'd654,  -14'd529,  14'd500,  -14'd118,  14'd1041,  14'd1484,  14'd1202,  -14'd470,  -14'd131,  14'd1251,  14'd96,  14'd1452,  
-14'd721,  14'd817,  14'd509,  -14'd591,  -14'd966,  -14'd1037,  -14'd1517,  -14'd779,  -14'd1558,  -14'd15,  -14'd392,  -14'd610,  -14'd996,  -14'd1031,  14'd789,  14'd1225,  
14'd590,  14'd1459,  -14'd367,  -14'd931,  14'd944,  14'd502,  14'd310,  -14'd577,  14'd1186,  -14'd1337,  -14'd905,  14'd1750,  -14'd1260,  -14'd505,  -14'd536,  -14'd606,  
14'd340,  -14'd1356,  -14'd245,  -14'd933,  14'd44,  -14'd491,  14'd1685,  -14'd1059,  -14'd122,  -14'd532,  -14'd333,  14'd133,  -14'd1235,  -14'd461,  14'd1207,  -14'd838,  
14'd1311,  -14'd79,  14'd508,  -14'd492,  14'd636,  -14'd1190,  14'd111,  -14'd457,  14'd144,  14'd524,  -14'd1069,  -14'd970,  -14'd1201,  14'd1363,  -14'd313,  -14'd265,  
-14'd432,  14'd19,  -14'd106,  -14'd109,  -14'd726,  14'd114,  -14'd789,  14'd693,  14'd615,  14'd31,  -14'd88,  -14'd2,  -14'd817,  14'd1896,  14'd1217,  -14'd173,  
14'd259,  -14'd1011,  14'd2327,  14'd1319,  14'd189,  14'd119,  14'd641,  14'd893,  -14'd367,  -14'd922,  -14'd859,  14'd309,  14'd1188,  -14'd532,  14'd2401,  14'd1359,  

14'd605,  -14'd14,  -14'd995,  -14'd1712,  -14'd1675,  14'd1528,  14'd1240,  14'd295,  14'd1601,  -14'd1095,  14'd386,  14'd395,  -14'd266,  14'd927,  -14'd933,  -14'd87,  
-14'd193,  -14'd1545,  -14'd962,  14'd464,  -14'd132,  14'd751,  -14'd951,  -14'd1422,  -14'd250,  -14'd1145,  14'd386,  -14'd36,  -14'd178,  -14'd549,  14'd1200,  14'd709,  
14'd889,  14'd210,  -14'd702,  14'd736,  -14'd1090,  14'd802,  -14'd495,  14'd443,  14'd329,  -14'd313,  14'd240,  -14'd1030,  -14'd473,  -14'd1175,  -14'd292,  -14'd49,  
-14'd1198,  -14'd6,  -14'd138,  14'd1147,  14'd817,  14'd529,  -14'd723,  -14'd911,  -14'd390,  14'd249,  14'd794,  -14'd449,  14'd862,  -14'd2955,  14'd409,  14'd741,  
-14'd1803,  -14'd1785,  14'd572,  14'd250,  14'd1010,  -14'd1207,  -14'd635,  14'd624,  -14'd356,  -14'd1010,  14'd704,  -14'd581,  14'd780,  14'd1083,  -14'd376,  14'd1933,  
14'd417,  14'd714,  -14'd265,  14'd1109,  -14'd70,  14'd584,  -14'd1366,  -14'd559,  -14'd1384,  14'd1965,  -14'd1592,  14'd15,  -14'd644,  -14'd540,  14'd37,  14'd504,  
14'd579,  -14'd225,  14'd391,  14'd1618,  -14'd1346,  -14'd51,  -14'd2311,  14'd1009,  14'd1082,  -14'd732,  -14'd327,  -14'd1352,  14'd1482,  14'd126,  14'd979,  14'd621,  
-14'd1330,  14'd164,  14'd33,  -14'd792,  -14'd719,  14'd129,  14'd362,  14'd100,  14'd1604,  14'd1734,  14'd2688,  -14'd557,  14'd271,  -14'd163,  -14'd551,  -14'd29,  
-14'd2818,  -14'd1315,  -14'd300,  -14'd774,  -14'd846,  -14'd519,  14'd812,  14'd954,  14'd295,  14'd2035,  14'd48,  -14'd234,  14'd278,  -14'd541,  14'd1052,  14'd403,  
-14'd993,  14'd8,  14'd414,  -14'd428,  -14'd1139,  14'd531,  -14'd717,  -14'd249,  14'd867,  14'd594,  14'd1057,  14'd730,  14'd623,  -14'd1677,  14'd220,  14'd685,  
14'd859,  14'd17,  -14'd860,  -14'd164,  14'd989,  -14'd368,  -14'd3204,  -14'd7,  14'd966,  14'd1130,  14'd715,  -14'd555,  14'd770,  -14'd106,  -14'd221,  -14'd34,  
-14'd640,  14'd1123,  14'd627,  -14'd1062,  14'd70,  14'd465,  -14'd955,  14'd1719,  14'd830,  14'd335,  -14'd845,  14'd873,  -14'd130,  14'd279,  -14'd215,  -14'd798,  
14'd805,  -14'd694,  -14'd1221,  14'd436,  14'd1382,  14'd488,  14'd232,  -14'd1099,  -14'd103,  -14'd617,  14'd534,  14'd642,  14'd1305,  -14'd741,  14'd701,  -14'd1159,  
-14'd666,  14'd1191,  14'd181,  -14'd659,  14'd491,  -14'd1145,  -14'd168,  14'd528,  -14'd717,  14'd636,  14'd1234,  -14'd215,  -14'd682,  -14'd168,  -14'd242,  -14'd403,  
14'd756,  14'd839,  -14'd426,  -14'd463,  14'd298,  14'd1277,  14'd770,  14'd381,  14'd186,  -14'd28,  14'd510,  -14'd682,  14'd1432,  -14'd545,  14'd482,  -14'd281,  
14'd642,  -14'd47,  14'd259,  14'd949,  14'd1732,  14'd274,  14'd1682,  -14'd800,  14'd1915,  14'd1228,  -14'd59,  -14'd444,  14'd424,  14'd915,  14'd726,  14'd1462,  
14'd1598,  14'd821,  14'd290,  14'd223,  -14'd445,  14'd264,  -14'd715,  -14'd338,  14'd414,  14'd728,  14'd747,  14'd1831,  14'd2004,  14'd201,  14'd388,  14'd953,  
-14'd331,  -14'd4,  -14'd169,  14'd1136,  14'd347,  -14'd907,  14'd179,  -14'd911,  14'd464,  14'd1509,  -14'd404,  -14'd887,  -14'd2,  -14'd1229,  -14'd626,  14'd459,  
-14'd452,  -14'd410,  -14'd943,  -14'd575,  14'd506,  -14'd834,  14'd114,  -14'd694,  -14'd166,  14'd4,  -14'd1044,  -14'd673,  -14'd1022,  -14'd694,  14'd855,  14'd1079,  
14'd960,  -14'd1348,  14'd1457,  14'd698,  -14'd361,  14'd1435,  14'd42,  -14'd445,  14'd560,  14'd2752,  14'd249,  -14'd1173,  14'd262,  14'd1095,  -14'd218,  14'd391,  
14'd155,  -14'd238,  -14'd273,  14'd1052,  14'd550,  14'd725,  14'd1174,  14'd1615,  14'd1233,  14'd982,  14'd768,  -14'd986,  14'd1318,  -14'd448,  -14'd58,  -14'd493,  
14'd889,  -14'd1932,  -14'd738,  -14'd986,  14'd943,  -14'd762,  -14'd538,  14'd222,  -14'd452,  -14'd330,  14'd98,  -14'd361,  14'd511,  14'd760,  -14'd99,  14'd217,  
-14'd1235,  -14'd849,  -14'd866,  -14'd282,  14'd150,  14'd102,  -14'd671,  -14'd996,  14'd197,  14'd197,  -14'd505,  14'd1697,  -14'd445,  14'd157,  14'd245,  -14'd176,  
14'd484,  -14'd275,  -14'd1022,  14'd386,  14'd568,  -14'd342,  -14'd624,  -14'd59,  14'd839,  -14'd891,  14'd223,  -14'd666,  -14'd524,  14'd705,  -14'd622,  14'd931,  
-14'd52,  14'd171,  14'd222,  14'd775,  -14'd4,  14'd724,  -14'd74,  14'd817,  -14'd317,  -14'd487,  14'd851,  -14'd150,  14'd193,  -14'd619,  14'd841,  14'd1428,  

-14'd891,  14'd487,  14'd977,  -14'd1021,  14'd966,  -14'd1641,  14'd385,  -14'd1850,  14'd652,  14'd530,  14'd625,  -14'd905,  14'd531,  14'd1847,  14'd391,  14'd1163,  
-14'd1378,  -14'd1310,  14'd1043,  -14'd85,  14'd133,  -14'd483,  14'd1332,  -14'd1417,  14'd99,  -14'd1077,  14'd453,  14'd355,  -14'd732,  14'd1926,  -14'd431,  14'd649,  
14'd1104,  -14'd629,  14'd1219,  -14'd894,  -14'd2315,  14'd129,  -14'd105,  -14'd495,  -14'd956,  -14'd630,  14'd1411,  -14'd1570,  -14'd1163,  14'd2460,  14'd576,  -14'd814,  
14'd919,  14'd573,  -14'd980,  -14'd1426,  -14'd672,  -14'd248,  14'd1064,  14'd1014,  14'd594,  -14'd273,  -14'd494,  14'd66,  14'd1219,  -14'd1216,  14'd920,  -14'd151,  
14'd522,  14'd3411,  -14'd1920,  14'd1231,  -14'd372,  14'd423,  14'd734,  -14'd129,  -14'd148,  14'd48,  14'd1705,  14'd354,  14'd2318,  14'd499,  14'd72,  14'd2118,  
-14'd1213,  -14'd373,  14'd755,  -14'd531,  -14'd1236,  -14'd1029,  14'd1067,  -14'd614,  -14'd804,  -14'd361,  14'd1505,  -14'd60,  14'd420,  14'd1086,  14'd463,  14'd536,  
14'd688,  14'd51,  -14'd381,  14'd579,  14'd957,  -14'd1023,  14'd1608,  14'd680,  -14'd23,  -14'd77,  14'd1586,  14'd460,  14'd60,  14'd786,  -14'd1336,  -14'd1225,  
14'd234,  -14'd1458,  14'd541,  -14'd1643,  14'd255,  14'd144,  -14'd496,  14'd68,  14'd2077,  -14'd57,  14'd300,  14'd258,  -14'd162,  -14'd615,  -14'd1283,  -14'd745,  
14'd827,  14'd2008,  14'd99,  14'd567,  14'd217,  -14'd17,  -14'd793,  14'd2430,  14'd637,  14'd548,  14'd1582,  -14'd249,  -14'd309,  -14'd582,  14'd374,  -14'd1135,  
14'd175,  14'd392,  14'd508,  -14'd32,  14'd863,  14'd1179,  -14'd117,  14'd1424,  -14'd70,  14'd2435,  14'd429,  14'd190,  -14'd314,  14'd829,  14'd1820,  14'd16,  
14'd1291,  14'd111,  14'd659,  -14'd699,  -14'd2859,  14'd1248,  14'd2106,  -14'd550,  -14'd1352,  14'd606,  14'd661,  14'd771,  -14'd320,  -14'd163,  14'd692,  14'd1691,  
-14'd487,  14'd695,  14'd953,  14'd145,  14'd630,  -14'd665,  14'd408,  14'd500,  14'd11,  14'd73,  -14'd819,  -14'd341,  -14'd368,  14'd1654,  -14'd189,  -14'd312,  
-14'd924,  14'd395,  14'd79,  -14'd959,  14'd705,  -14'd886,  -14'd564,  -14'd347,  -14'd491,  -14'd562,  -14'd10,  -14'd202,  14'd914,  -14'd340,  -14'd1011,  14'd422,  
-14'd782,  -14'd735,  -14'd1546,  -14'd327,  14'd395,  -14'd609,  -14'd1739,  -14'd1107,  -14'd716,  14'd1423,  -14'd755,  14'd316,  -14'd354,  -14'd1499,  14'd979,  14'd1305,  
-14'd389,  14'd165,  14'd749,  -14'd20,  14'd934,  -14'd308,  -14'd1308,  -14'd685,  14'd495,  14'd255,  14'd572,  14'd615,  -14'd91,  -14'd562,  14'd1887,  14'd786,  
14'd171,  14'd445,  14'd1658,  14'd177,  -14'd723,  14'd453,  -14'd220,  14'd2251,  14'd209,  14'd62,  14'd391,  -14'd5,  -14'd54,  14'd82,  14'd766,  14'd259,  
-14'd498,  14'd758,  14'd407,  14'd1640,  -14'd1053,  14'd374,  -14'd122,  14'd13,  -14'd1792,  -14'd854,  -14'd409,  -14'd1396,  -14'd1250,  14'd343,  14'd459,  -14'd1521,  
14'd612,  -14'd1085,  14'd647,  14'd550,  14'd1152,  -14'd722,  14'd5,  14'd345,  14'd863,  -14'd1188,  -14'd52,  -14'd196,  14'd1058,  14'd1035,  -14'd701,  -14'd1293,  
14'd170,  -14'd289,  -14'd1285,  -14'd366,  14'd1581,  14'd1146,  14'd138,  -14'd171,  14'd250,  14'd6,  14'd1404,  14'd490,  14'd12,  14'd21,  -14'd123,  14'd54,  
14'd1085,  14'd1920,  14'd1728,  -14'd1103,  14'd350,  14'd248,  14'd751,  14'd145,  14'd292,  -14'd470,  -14'd66,  14'd1020,  14'd356,  -14'd533,  14'd512,  -14'd11,  
-14'd1717,  -14'd148,  -14'd159,  -14'd213,  -14'd456,  14'd892,  -14'd345,  14'd176,  14'd133,  -14'd79,  -14'd597,  14'd779,  -14'd910,  14'd470,  -14'd686,  14'd156,  
-14'd1673,  -14'd613,  14'd363,  14'd1037,  14'd778,  14'd1721,  14'd1467,  14'd83,  14'd1066,  -14'd252,  14'd810,  -14'd267,  14'd1390,  -14'd530,  -14'd239,  14'd91,  
-14'd988,  14'd221,  -14'd538,  14'd203,  14'd271,  14'd1067,  14'd403,  14'd389,  14'd1456,  -14'd376,  14'd1580,  14'd241,  -14'd336,  -14'd675,  -14'd847,  14'd960,  
14'd1884,  14'd207,  14'd1754,  14'd352,  -14'd96,  -14'd515,  -14'd1198,  14'd1234,  -14'd157,  14'd500,  14'd970,  14'd982,  14'd564,  14'd317,  -14'd1818,  -14'd877,  
14'd1394,  14'd78,  14'd1032,  -14'd147,  14'd680,  -14'd273,  14'd758,  -14'd474,  14'd1555,  14'd684,  -14'd622,  14'd2298,  14'd748,  -14'd1376,  14'd11,  -14'd255,  

-14'd1631,  -14'd217,  -14'd835,  14'd158,  14'd535,  14'd171,  -14'd1346,  14'd1256,  -14'd843,  14'd277,  -14'd269,  -14'd1400,  14'd2190,  -14'd298,  -14'd261,  -14'd1424,  
-14'd507,  14'd747,  14'd127,  -14'd54,  14'd798,  14'd919,  -14'd759,  14'd36,  14'd508,  14'd448,  -14'd1360,  -14'd261,  14'd725,  -14'd273,  14'd834,  14'd166,  
-14'd1071,  -14'd283,  14'd1717,  14'd226,  -14'd1399,  14'd714,  14'd673,  -14'd1171,  14'd98,  -14'd784,  14'd273,  -14'd787,  -14'd590,  14'd1346,  14'd991,  14'd1593,  
-14'd375,  -14'd748,  14'd89,  14'd1819,  -14'd1590,  -14'd1162,  -14'd810,  -14'd22,  14'd1789,  14'd439,  14'd1089,  14'd40,  -14'd1098,  14'd169,  14'd235,  -14'd468,  
-14'd39,  -14'd1120,  14'd781,  -14'd540,  14'd1467,  -14'd1051,  -14'd877,  -14'd949,  -14'd317,  -14'd571,  14'd1127,  14'd213,  -14'd349,  14'd213,  -14'd167,  14'd122,  
-14'd1329,  -14'd404,  -14'd1913,  14'd1110,  14'd759,  -14'd1556,  -14'd350,  -14'd1596,  14'd240,  -14'd1072,  14'd1005,  -14'd471,  14'd480,  -14'd71,  -14'd1277,  14'd617,  
-14'd879,  -14'd980,  -14'd1686,  14'd957,  14'd1987,  -14'd829,  -14'd806,  -14'd346,  -14'd570,  14'd746,  -14'd803,  14'd1146,  14'd1357,  -14'd796,  -14'd51,  14'd919,  
-14'd216,  14'd284,  14'd191,  14'd590,  14'd378,  -14'd412,  -14'd27,  -14'd152,  -14'd669,  14'd24,  14'd751,  14'd520,  14'd986,  -14'd224,  -14'd1963,  -14'd103,  
-14'd100,  14'd120,  14'd420,  -14'd861,  -14'd458,  14'd974,  -14'd824,  -14'd802,  -14'd735,  14'd740,  14'd861,  14'd168,  14'd456,  14'd1769,  -14'd45,  -14'd156,  
14'd556,  14'd1710,  14'd1333,  14'd876,  -14'd389,  -14'd1086,  14'd1019,  -14'd95,  14'd853,  14'd798,  14'd212,  14'd16,  -14'd1008,  14'd1047,  14'd1761,  -14'd573,  
-14'd789,  14'd535,  -14'd1234,  -14'd1420,  -14'd917,  14'd1144,  -14'd1850,  14'd511,  14'd1441,  -14'd871,  14'd1612,  14'd452,  -14'd185,  -14'd81,  14'd868,  14'd868,  
14'd883,  14'd178,  14'd31,  14'd356,  14'd432,  14'd848,  -14'd734,  -14'd1291,  14'd451,  14'd2242,  14'd207,  14'd224,  14'd543,  -14'd1340,  -14'd1196,  14'd1903,  
14'd638,  14'd546,  -14'd1565,  14'd522,  14'd1850,  -14'd1419,  14'd166,  14'd624,  -14'd675,  14'd666,  14'd1296,  14'd1225,  14'd132,  -14'd519,  14'd19,  14'd1595,  
14'd270,  14'd773,  14'd745,  14'd348,  14'd799,  -14'd469,  14'd735,  14'd656,  14'd1174,  14'd1198,  14'd1142,  -14'd532,  -14'd941,  14'd167,  -14'd1368,  -14'd1755,  
14'd1004,  14'd439,  14'd172,  14'd832,  -14'd1585,  14'd976,  14'd347,  -14'd276,  14'd459,  -14'd1023,  -14'd1196,  -14'd171,  14'd1279,  -14'd895,  -14'd2017,  -14'd182,  
14'd72,  -14'd321,  -14'd987,  -14'd162,  -14'd1500,  -14'd538,  -14'd1048,  -14'd528,  14'd663,  -14'd65,  14'd1502,  -14'd490,  -14'd313,  -14'd1219,  14'd121,  14'd741,  
-14'd927,  14'd45,  -14'd1326,  14'd637,  14'd550,  -14'd49,  -14'd968,  14'd1489,  -14'd499,  14'd259,  14'd802,  14'd1012,  14'd465,  -14'd697,  14'd429,  14'd1010,  
14'd721,  14'd1245,  -14'd1467,  14'd425,  14'd731,  14'd303,  -14'd275,  14'd277,  14'd326,  -14'd936,  14'd815,  14'd1052,  14'd591,  14'd837,  -14'd616,  -14'd273,  
14'd393,  -14'd440,  -14'd1376,  14'd1760,  14'd294,  -14'd793,  -14'd181,  14'd89,  14'd393,  -14'd814,  14'd1576,  -14'd597,  14'd1007,  -14'd28,  14'd212,  14'd933,  
14'd828,  -14'd690,  -14'd1259,  14'd676,  14'd1360,  14'd1210,  -14'd241,  -14'd717,  14'd962,  -14'd134,  14'd154,  14'd86,  14'd2462,  14'd250,  -14'd118,  14'd242,  
-14'd159,  -14'd683,  -14'd347,  -14'd1016,  -14'd294,  -14'd33,  14'd1497,  -14'd1448,  -14'd1370,  14'd1064,  14'd571,  -14'd588,  14'd877,  14'd36,  14'd721,  14'd860,  
-14'd102,  14'd1535,  14'd575,  -14'd436,  14'd123,  -14'd1825,  -14'd308,  -14'd5,  -14'd37,  -14'd514,  14'd1371,  -14'd645,  14'd7,  -14'd2054,  14'd227,  14'd584,  
14'd843,  14'd562,  -14'd739,  -14'd72,  14'd1034,  -14'd341,  -14'd508,  -14'd681,  -14'd821,  14'd2057,  -14'd729,  -14'd54,  14'd696,  -14'd381,  14'd771,  -14'd943,  
-14'd1250,  14'd1810,  -14'd172,  14'd648,  14'd63,  -14'd993,  -14'd478,  -14'd101,  -14'd101,  14'd153,  14'd112,  -14'd1623,  14'd1513,  14'd253,  -14'd521,  -14'd1011,  
14'd188,  14'd1341,  14'd458,  -14'd630,  -14'd228,  14'd902,  -14'd1860,  14'd854,  14'd398,  14'd1329,  -14'd1345,  14'd503,  -14'd640,  -14'd653,  14'd239,  -14'd435,  

14'd428,  14'd7,  -14'd963,  -14'd108,  -14'd128,  14'd232,  14'd12,  -14'd467,  14'd1036,  -14'd463,  -14'd602,  14'd555,  14'd817,  -14'd254,  -14'd1116,  14'd633,  
14'd1119,  -14'd442,  14'd500,  14'd635,  -14'd1088,  14'd506,  -14'd125,  14'd92,  -14'd1503,  14'd690,  -14'd1206,  -14'd35,  -14'd1211,  -14'd1002,  -14'd1375,  -14'd733,  
-14'd459,  -14'd943,  -14'd299,  -14'd97,  14'd129,  14'd163,  -14'd32,  -14'd748,  14'd513,  -14'd692,  -14'd217,  -14'd915,  -14'd558,  -14'd506,  -14'd553,  14'd505,  
-14'd852,  -14'd564,  -14'd730,  14'd3,  -14'd63,  -14'd208,  14'd262,  14'd495,  14'd392,  -14'd720,  -14'd286,  14'd616,  -14'd547,  -14'd1313,  -14'd127,  -14'd566,  
14'd129,  14'd675,  14'd757,  -14'd743,  -14'd212,  -14'd740,  -14'd235,  14'd12,  14'd420,  14'd31,  -14'd1199,  -14'd54,  14'd98,  14'd488,  14'd1088,  14'd610,  
-14'd478,  -14'd524,  -14'd472,  -14'd649,  14'd157,  14'd537,  -14'd936,  -14'd846,  14'd25,  -14'd1442,  14'd717,  14'd128,  -14'd710,  14'd705,  -14'd401,  -14'd369,  
14'd974,  14'd11,  14'd596,  -14'd782,  14'd667,  -14'd982,  -14'd70,  -14'd683,  -14'd547,  -14'd630,  14'd528,  14'd45,  14'd1007,  -14'd276,  14'd314,  14'd543,  
14'd140,  -14'd870,  -14'd687,  -14'd384,  14'd480,  -14'd201,  -14'd1695,  14'd812,  -14'd366,  14'd37,  14'd349,  -14'd1309,  14'd1010,  -14'd209,  -14'd231,  -14'd1061,  
14'd1200,  -14'd451,  14'd47,  -14'd40,  14'd170,  14'd1327,  -14'd1109,  14'd450,  -14'd974,  -14'd750,  -14'd387,  14'd296,  14'd868,  -14'd644,  14'd881,  14'd531,  
14'd1028,  -14'd208,  14'd560,  14'd1452,  -14'd141,  -14'd662,  -14'd1424,  14'd1167,  14'd163,  -14'd1473,  -14'd372,  -14'd150,  -14'd214,  -14'd90,  14'd935,  14'd927,  
-14'd110,  14'd128,  -14'd271,  -14'd546,  -14'd1440,  14'd293,  -14'd766,  -14'd367,  -14'd714,  -14'd1530,  -14'd312,  14'd71,  14'd226,  -14'd169,  14'd806,  -14'd1340,  
14'd998,  -14'd363,  14'd980,  14'd657,  -14'd1703,  14'd713,  -14'd315,  14'd371,  -14'd1432,  14'd1315,  14'd692,  14'd73,  14'd620,  -14'd767,  14'd87,  14'd178,  
14'd14,  -14'd684,  -14'd1127,  -14'd98,  14'd49,  -14'd1476,  14'd240,  -14'd317,  14'd684,  14'd302,  -14'd519,  14'd365,  -14'd253,  14'd178,  14'd618,  14'd505,  
-14'd464,  14'd518,  -14'd757,  -14'd15,  -14'd56,  -14'd717,  -14'd657,  -14'd877,  -14'd1471,  -14'd1457,  -14'd708,  -14'd782,  -14'd819,  14'd239,  -14'd677,  -14'd271,  
-14'd953,  14'd69,  -14'd1082,  -14'd746,  -14'd601,  -14'd218,  -14'd79,  -14'd1391,  -14'd64,  -14'd645,  -14'd1267,  -14'd323,  14'd28,  -14'd154,  14'd590,  14'd71,  
-14'd402,  -14'd27,  -14'd150,  -14'd101,  14'd318,  -14'd565,  -14'd521,  14'd175,  14'd879,  -14'd501,  -14'd711,  -14'd442,  -14'd633,  -14'd260,  14'd626,  14'd990,  
14'd668,  14'd1230,  14'd542,  -14'd861,  -14'd181,  14'd948,  -14'd1519,  -14'd41,  14'd261,  -14'd363,  14'd324,  14'd138,  -14'd88,  14'd410,  -14'd765,  14'd684,  
-14'd1459,  14'd62,  -14'd154,  14'd159,  -14'd1078,  14'd1000,  14'd584,  -14'd27,  -14'd1193,  -14'd871,  -14'd3,  -14'd563,  -14'd1057,  -14'd495,  14'd363,  -14'd123,  
14'd1060,  -14'd102,  -14'd668,  14'd753,  14'd1061,  14'd580,  -14'd107,  -14'd730,  14'd945,  -14'd388,  -14'd581,  14'd122,  14'd1349,  14'd248,  14'd413,  -14'd71,  
14'd1196,  -14'd1291,  -14'd531,  -14'd771,  -14'd386,  -14'd461,  -14'd686,  -14'd84,  -14'd827,  14'd710,  14'd178,  14'd149,  -14'd313,  14'd1100,  -14'd552,  14'd713,  
-14'd297,  14'd496,  -14'd24,  14'd1153,  -14'd1486,  14'd614,  14'd382,  -14'd310,  14'd132,  -14'd1200,  -14'd149,  -14'd972,  14'd566,  -14'd1103,  -14'd1202,  -14'd1475,  
-14'd419,  14'd93,  -14'd634,  14'd1195,  14'd372,  -14'd1533,  -14'd225,  -14'd684,  14'd384,  14'd761,  14'd443,  14'd491,  -14'd1689,  -14'd445,  -14'd543,  -14'd1003,  
-14'd286,  14'd51,  -14'd1210,  -14'd647,  14'd220,  14'd298,  -14'd785,  -14'd735,  14'd126,  -14'd1210,  14'd1146,  -14'd1436,  -14'd476,  -14'd1225,  14'd809,  -14'd1065,  
-14'd744,  -14'd487,  14'd268,  -14'd353,  -14'd767,  14'd1413,  -14'd106,  -14'd468,  -14'd262,  14'd913,  -14'd718,  14'd653,  -14'd928,  -14'd344,  14'd300,  -14'd862,  
14'd195,  14'd338,  14'd53,  -14'd231,  14'd353,  -14'd820,  14'd8,  -14'd909,  14'd1290,  -14'd772,  14'd1031,  -14'd699,  -14'd1289,  -14'd157,  14'd109,  -14'd511,  

-14'd887,  -14'd129,  -14'd616,  -14'd21,  14'd363,  14'd865,  14'd332,  -14'd949,  -14'd1636,  14'd4,  -14'd303,  14'd845,  -14'd499,  -14'd826,  -14'd1064,  -14'd712,  
14'd112,  -14'd339,  -14'd1479,  -14'd90,  -14'd496,  14'd301,  -14'd284,  14'd422,  -14'd67,  14'd310,  14'd384,  14'd740,  -14'd1014,  -14'd1996,  -14'd444,  14'd316,  
-14'd1712,  -14'd828,  -14'd523,  -14'd388,  14'd2086,  14'd527,  -14'd800,  -14'd987,  -14'd1275,  14'd642,  14'd281,  -14'd81,  14'd1644,  -14'd3233,  -14'd266,  -14'd27,  
-14'd1948,  -14'd1670,  14'd655,  14'd472,  14'd113,  -14'd1588,  -14'd147,  14'd263,  -14'd1008,  -14'd20,  -14'd427,  14'd741,  14'd237,  -14'd37,  14'd376,  -14'd560,  
-14'd369,  -14'd465,  -14'd173,  -14'd888,  14'd1435,  -14'd577,  -14'd651,  14'd1094,  14'd715,  -14'd588,  14'd278,  14'd576,  -14'd620,  -14'd378,  -14'd391,  -14'd166,  
-14'd1470,  14'd615,  14'd84,  -14'd847,  -14'd1082,  -14'd1427,  -14'd7,  14'd752,  14'd1390,  -14'd640,  14'd1914,  14'd670,  14'd479,  14'd435,  14'd214,  14'd269,  
14'd183,  14'd973,  14'd822,  14'd136,  14'd172,  -14'd1228,  14'd592,  -14'd972,  -14'd54,  14'd1179,  -14'd1431,  14'd845,  14'd899,  -14'd862,  14'd1438,  14'd871,  
-14'd851,  -14'd883,  -14'd1450,  -14'd30,  14'd676,  -14'd542,  14'd152,  -14'd766,  -14'd388,  -14'd352,  14'd199,  14'd1284,  14'd1067,  -14'd2200,  14'd1118,  -14'd27,  
14'd504,  -14'd368,  -14'd415,  14'd352,  -14'd342,  -14'd159,  14'd825,  14'd776,  14'd967,  14'd143,  14'd170,  14'd501,  14'd1111,  14'd991,  14'd595,  14'd1570,  
14'd927,  14'd678,  14'd410,  14'd1714,  14'd92,  14'd738,  14'd170,  14'd528,  -14'd714,  -14'd1841,  -14'd90,  -14'd45,  14'd323,  14'd612,  -14'd679,  -14'd25,  
14'd235,  14'd102,  -14'd890,  -14'd360,  14'd542,  -14'd228,  -14'd1947,  14'd99,  14'd727,  14'd571,  -14'd1530,  -14'd695,  14'd1474,  14'd750,  14'd668,  14'd537,  
-14'd45,  14'd594,  -14'd875,  14'd260,  -14'd173,  -14'd834,  -14'd1469,  -14'd329,  -14'd1196,  14'd471,  14'd1282,  -14'd1174,  -14'd101,  14'd889,  14'd646,  -14'd68,  
14'd1089,  -14'd1372,  14'd411,  14'd1172,  -14'd887,  14'd589,  -14'd1006,  -14'd56,  -14'd1219,  14'd460,  14'd506,  14'd1540,  -14'd237,  -14'd2504,  14'd77,  -14'd445,  
14'd827,  -14'd1837,  -14'd379,  -14'd151,  14'd1390,  -14'd732,  14'd578,  -14'd810,  14'd42,  14'd1351,  -14'd681,  14'd363,  14'd661,  14'd196,  14'd184,  14'd969,  
-14'd583,  -14'd850,  -14'd364,  -14'd1075,  14'd1143,  -14'd184,  14'd924,  -14'd1887,  -14'd690,  14'd600,  14'd583,  -14'd1072,  -14'd77,  -14'd59,  14'd237,  14'd1853,  
-14'd1627,  -14'd527,  -14'd1611,  -14'd584,  14'd1061,  -14'd1457,  -14'd1267,  -14'd666,  -14'd215,  -14'd161,  -14'd590,  -14'd444,  -14'd909,  -14'd925,  -14'd814,  14'd546,  
14'd1223,  14'd538,  -14'd297,  14'd1273,  14'd2090,  -14'd818,  -14'd1092,  -14'd1188,  14'd1253,  14'd728,  -14'd981,  14'd144,  14'd139,  -14'd1858,  -14'd506,  14'd292,  
-14'd384,  14'd767,  14'd768,  14'd813,  -14'd1235,  14'd919,  -14'd410,  14'd1037,  14'd237,  -14'd376,  14'd317,  -14'd206,  -14'd553,  -14'd2615,  14'd1027,  -14'd240,  
14'd379,  14'd940,  -14'd438,  -14'd319,  -14'd185,  -14'd376,  14'd521,  14'd458,  14'd1701,  -14'd693,  -14'd59,  14'd549,  14'd462,  14'd1125,  -14'd467,  -14'd506,  
-14'd108,  14'd169,  -14'd386,  -14'd282,  -14'd1711,  -14'd918,  14'd1066,  -14'd1745,  14'd1132,  -14'd521,  14'd528,  -14'd1661,  -14'd914,  -14'd724,  -14'd994,  -14'd739,  
14'd482,  -14'd209,  -14'd685,  -14'd1444,  -14'd705,  -14'd205,  14'd795,  -14'd715,  14'd1910,  -14'd91,  14'd1548,  14'd895,  14'd992,  -14'd1565,  14'd716,  14'd106,  
14'd1678,  -14'd1036,  -14'd394,  -14'd75,  14'd482,  14'd242,  -14'd204,  14'd496,  14'd981,  14'd757,  14'd432,  14'd985,  -14'd401,  -14'd203,  -14'd997,  -14'd113,  
14'd311,  14'd755,  14'd1089,  -14'd85,  -14'd1537,  -14'd118,  14'd895,  14'd1091,  14'd1548,  14'd1787,  14'd536,  14'd782,  14'd1169,  14'd720,  14'd193,  -14'd438,  
14'd394,  -14'd508,  14'd801,  -14'd244,  -14'd779,  -14'd765,  14'd466,  -14'd141,  -14'd533,  -14'd913,  14'd251,  14'd970,  14'd466,  14'd1602,  -14'd1056,  14'd1020,  
-14'd67,  -14'd949,  14'd920,  -14'd514,  -14'd1291,  14'd187,  14'd308,  -14'd134,  14'd1350,  -14'd444,  14'd6,  -14'd343,  -14'd154,  14'd508,  -14'd214,  -14'd749,  

14'd988,  -14'd943,  -14'd238,  -14'd1672,  -14'd318,  -14'd298,  -14'd1199,  14'd22,  14'd833,  14'd1035,  -14'd86,  -14'd373,  -14'd89,  14'd12,  14'd428,  14'd139,  
14'd1231,  -14'd273,  14'd371,  -14'd638,  14'd1029,  14'd170,  -14'd694,  -14'd884,  14'd798,  -14'd1691,  -14'd404,  -14'd1261,  -14'd1320,  -14'd276,  -14'd295,  14'd711,  
-14'd967,  -14'd476,  -14'd211,  14'd1183,  -14'd531,  14'd716,  14'd1133,  14'd1242,  -14'd1669,  -14'd1150,  -14'd689,  -14'd708,  -14'd1182,  14'd694,  14'd113,  14'd412,  
14'd258,  14'd842,  14'd452,  -14'd473,  14'd391,  -14'd111,  14'd1147,  -14'd540,  -14'd590,  14'd151,  14'd525,  -14'd291,  14'd1232,  -14'd572,  14'd191,  -14'd531,  
-14'd264,  14'd921,  14'd380,  -14'd991,  -14'd1070,  14'd1083,  -14'd297,  -14'd104,  -14'd754,  14'd353,  14'd123,  -14'd1176,  14'd176,  -14'd101,  -14'd1123,  14'd866,  
-14'd408,  14'd16,  -14'd601,  -14'd397,  -14'd663,  -14'd1074,  -14'd1072,  -14'd326,  14'd497,  -14'd958,  -14'd1058,  -14'd38,  14'd1188,  -14'd628,  -14'd819,  -14'd783,  
14'd390,  -14'd708,  14'd1418,  14'd1154,  -14'd450,  -14'd195,  -14'd804,  -14'd1296,  14'd987,  -14'd1,  -14'd590,  14'd261,  14'd43,  14'd111,  -14'd1301,  -14'd1694,  
-14'd279,  14'd647,  14'd353,  14'd191,  14'd522,  -14'd291,  -14'd721,  -14'd437,  -14'd1150,  -14'd212,  -14'd180,  14'd784,  14'd1137,  14'd362,  -14'd809,  -14'd440,  
14'd738,  -14'd636,  -14'd439,  -14'd719,  14'd1403,  14'd1101,  -14'd707,  -14'd1114,  -14'd770,  -14'd1389,  14'd701,  -14'd713,  14'd96,  14'd343,  -14'd724,  -14'd293,  
-14'd801,  -14'd764,  14'd939,  -14'd966,  14'd797,  -14'd296,  14'd1046,  -14'd969,  14'd375,  -14'd99,  -14'd216,  -14'd672,  -14'd1236,  14'd520,  -14'd920,  14'd582,  
-14'd920,  -14'd1019,  14'd341,  14'd588,  14'd112,  -14'd229,  -14'd329,  -14'd365,  -14'd180,  -14'd909,  -14'd1786,  -14'd1066,  14'd623,  14'd921,  14'd667,  -14'd157,  
14'd600,  14'd911,  -14'd658,  -14'd529,  -14'd368,  14'd47,  14'd832,  -14'd274,  -14'd236,  -14'd1166,  14'd309,  14'd450,  14'd385,  -14'd791,  -14'd1567,  14'd28,  
14'd231,  -14'd1208,  14'd9,  -14'd634,  -14'd298,  -14'd699,  14'd448,  -14'd898,  14'd314,  14'd80,  -14'd41,  -14'd307,  -14'd942,  -14'd280,  -14'd302,  14'd1218,  
-14'd738,  -14'd1314,  14'd137,  -14'd91,  14'd521,  -14'd781,  -14'd170,  -14'd978,  -14'd1498,  -14'd450,  -14'd817,  14'd201,  -14'd1196,  -14'd262,  14'd28,  14'd379,  
-14'd465,  -14'd539,  -14'd71,  -14'd388,  14'd210,  14'd19,  14'd759,  14'd30,  14'd1294,  -14'd47,  14'd464,  -14'd758,  -14'd37,  14'd328,  14'd1274,  -14'd374,  
14'd434,  14'd828,  14'd752,  14'd610,  -14'd1166,  14'd978,  14'd1452,  -14'd530,  14'd1020,  -14'd368,  -14'd529,  -14'd616,  14'd546,  -14'd1439,  14'd24,  -14'd1405,  
14'd476,  -14'd42,  -14'd871,  14'd272,  -14'd322,  -14'd731,  14'd143,  14'd1103,  -14'd109,  14'd832,  14'd1182,  -14'd1305,  14'd768,  -14'd1257,  14'd771,  14'd597,  
-14'd234,  -14'd1126,  -14'd1668,  14'd1010,  14'd287,  -14'd484,  14'd645,  -14'd1109,  14'd730,  14'd603,  -14'd322,  14'd212,  -14'd750,  14'd234,  -14'd441,  -14'd43,  
-14'd1486,  -14'd416,  -14'd224,  14'd89,  14'd24,  -14'd606,  -14'd468,  14'd79,  -14'd274,  -14'd325,  14'd347,  14'd1333,  -14'd1087,  -14'd66,  14'd11,  14'd53,  
-14'd1448,  14'd569,  14'd1177,  -14'd799,  -14'd871,  14'd53,  -14'd1085,  14'd883,  -14'd1376,  14'd56,  14'd790,  -14'd220,  14'd310,  -14'd254,  14'd530,  -14'd680,  
-14'd105,  -14'd1410,  -14'd1012,  -14'd15,  -14'd416,  -14'd601,  -14'd859,  -14'd1366,  14'd566,  -14'd233,  -14'd113,  -14'd541,  -14'd1206,  14'd717,  -14'd445,  -14'd83,  
14'd421,  14'd1098,  14'd198,  -14'd79,  14'd445,  -14'd153,  14'd196,  -14'd353,  14'd1317,  -14'd23,  14'd728,  14'd510,  -14'd9,  14'd506,  14'd219,  -14'd1,  
14'd891,  -14'd413,  -14'd108,  -14'd1540,  14'd284,  -14'd441,  14'd873,  -14'd450,  14'd41,  14'd416,  -14'd1085,  -14'd554,  -14'd17,  14'd242,  -14'd358,  -14'd1394,  
14'd313,  -14'd156,  14'd475,  -14'd611,  14'd56,  -14'd836,  14'd1300,  -14'd751,  -14'd368,  -14'd16,  14'd337,  -14'd258,  -14'd934,  -14'd387,  -14'd696,  -14'd474,  
14'd1104,  14'd295,  14'd489,  -14'd235,  -14'd625,  14'd550,  14'd767,  14'd200,  14'd220,  -14'd909,  14'd853,  -14'd367,  14'd252,  -14'd405,  -14'd989,  -14'd718,  

14'd237,  -14'd636,  14'd665,  -14'd599,  -14'd978,  -14'd160,  -14'd771,  -14'd248,  -14'd639,  14'd1053,  14'd634,  -14'd29,  14'd793,  -14'd319,  -14'd769,  -14'd1549,  
-14'd416,  14'd639,  -14'd926,  -14'd896,  -14'd1200,  14'd749,  14'd658,  -14'd1489,  14'd36,  -14'd895,  -14'd383,  -14'd597,  14'd98,  -14'd165,  14'd213,  14'd421,  
-14'd39,  14'd1453,  14'd280,  -14'd442,  -14'd9,  14'd784,  14'd167,  -14'd819,  14'd1087,  14'd1215,  14'd16,  -14'd512,  -14'd1301,  -14'd547,  -14'd814,  14'd88,  
14'd277,  -14'd1270,  -14'd1113,  14'd1120,  14'd871,  14'd1255,  14'd659,  -14'd1060,  -14'd465,  14'd624,  -14'd1178,  14'd505,  -14'd605,  -14'd1507,  -14'd1370,  -14'd527,  
14'd790,  -14'd243,  -14'd270,  -14'd935,  14'd1148,  14'd367,  14'd124,  -14'd474,  14'd398,  14'd646,  -14'd232,  -14'd258,  -14'd1289,  -14'd41,  14'd746,  14'd336,  
-14'd1029,  14'd1106,  -14'd1399,  -14'd1352,  -14'd1842,  14'd72,  -14'd68,  -14'd1270,  14'd615,  -14'd1329,  -14'd1285,  -14'd709,  -14'd794,  14'd350,  -14'd285,  -14'd280,  
-14'd1030,  -14'd524,  -14'd1005,  14'd805,  -14'd325,  -14'd1455,  -14'd1122,  -14'd614,  -14'd556,  -14'd1852,  -14'd998,  -14'd1039,  -14'd845,  -14'd551,  -14'd388,  -14'd931,  
-14'd658,  -14'd15,  -14'd1323,  -14'd849,  -14'd387,  -14'd620,  14'd891,  -14'd704,  -14'd1195,  14'd1355,  -14'd813,  -14'd511,  14'd73,  -14'd1750,  -14'd942,  14'd546,  
-14'd63,  -14'd810,  14'd178,  -14'd1205,  -14'd1073,  -14'd860,  -14'd48,  -14'd989,  14'd525,  -14'd295,  -14'd693,  14'd90,  14'd74,  -14'd899,  14'd113,  -14'd158,  
14'd11,  -14'd1619,  14'd915,  -14'd611,  14'd735,  14'd595,  14'd1024,  -14'd232,  14'd139,  14'd530,  -14'd631,  -14'd50,  14'd427,  -14'd254,  14'd948,  14'd170,  
-14'd1354,  14'd633,  -14'd251,  -14'd1171,  -14'd630,  -14'd832,  -14'd860,  14'd691,  14'd490,  14'd1001,  -14'd652,  -14'd932,  -14'd181,  14'd274,  14'd1034,  -14'd269,  
-14'd770,  -14'd500,  -14'd1228,  -14'd226,  -14'd11,  14'd288,  -14'd512,  -14'd1896,  14'd584,  -14'd428,  -14'd496,  14'd384,  -14'd544,  -14'd991,  14'd6,  -14'd194,  
14'd299,  -14'd1355,  -14'd668,  14'd502,  14'd715,  14'd240,  14'd290,  -14'd265,  -14'd1682,  -14'd693,  14'd310,  -14'd128,  -14'd615,  14'd229,  -14'd663,  14'd131,  
14'd263,  -14'd352,  -14'd1886,  14'd42,  14'd402,  -14'd338,  14'd41,  14'd169,  -14'd159,  14'd354,  14'd284,  -14'd457,  -14'd624,  14'd1032,  14'd143,  14'd196,  
-14'd447,  -14'd162,  -14'd337,  -14'd323,  14'd434,  -14'd624,  -14'd183,  -14'd943,  14'd61,  -14'd989,  -14'd1339,  14'd670,  14'd868,  14'd492,  -14'd789,  14'd169,  
-14'd1139,  14'd243,  -14'd28,  -14'd1117,  14'd9,  -14'd331,  14'd44,  -14'd1120,  -14'd478,  -14'd417,  -14'd114,  -14'd750,  -14'd421,  14'd294,  -14'd378,  14'd551,  
-14'd2,  -14'd29,  -14'd38,  -14'd320,  14'd79,  -14'd1216,  -14'd107,  14'd226,  -14'd1345,  14'd804,  14'd42,  -14'd1334,  -14'd1238,  14'd750,  14'd1214,  14'd522,  
-14'd1294,  -14'd623,  14'd426,  -14'd395,  -14'd287,  -14'd1124,  -14'd354,  14'd925,  14'd1587,  14'd520,  -14'd1587,  -14'd871,  -14'd620,  14'd154,  14'd243,  -14'd626,  
-14'd805,  14'd947,  -14'd1985,  -14'd675,  -14'd649,  -14'd233,  14'd90,  -14'd419,  -14'd1236,  -14'd774,  -14'd1361,  14'd395,  -14'd68,  -14'd487,  -14'd1170,  -14'd210,  
14'd179,  -14'd1332,  -14'd412,  -14'd1136,  -14'd83,  -14'd631,  -14'd533,  -14'd1219,  -14'd206,  -14'd296,  -14'd840,  -14'd1402,  14'd200,  -14'd47,  14'd319,  14'd691,  
-14'd825,  -14'd33,  -14'd686,  -14'd1820,  -14'd410,  -14'd338,  14'd356,  14'd411,  14'd416,  -14'd1523,  -14'd227,  -14'd405,  14'd242,  -14'd33,  14'd169,  -14'd450,  
14'd850,  -14'd450,  -14'd859,  -14'd965,  -14'd553,  14'd714,  14'd561,  -14'd1299,  14'd669,  14'd197,  14'd381,  14'd66,  14'd161,  14'd479,  14'd17,  -14'd991,  
14'd454,  -14'd452,  -14'd1323,  14'd813,  14'd690,  14'd595,  14'd233,  -14'd830,  -14'd421,  14'd217,  14'd1180,  14'd87,  -14'd82,  -14'd1097,  14'd1,  14'd640,  
14'd768,  -14'd994,  -14'd637,  -14'd372,  -14'd655,  -14'd1032,  -14'd677,  -14'd536,  14'd674,  -14'd1005,  -14'd264,  -14'd11,  -14'd60,  14'd45,  14'd106,  14'd238,  
-14'd299,  14'd564,  -14'd289,  -14'd366,  14'd490,  -14'd712,  -14'd1265,  -14'd823,  14'd183,  -14'd1388,  14'd1044,  -14'd585,  -14'd1248,  -14'd586,  14'd398,  14'd512,  

14'd788,  14'd1011,  14'd2234,  14'd1337,  -14'd190,  14'd99,  -14'd1472,  14'd92,  -14'd379,  14'd825,  -14'd396,  -14'd145,  14'd965,  14'd731,  14'd1289,  -14'd744,  
14'd1063,  14'd626,  -14'd653,  -14'd40,  14'd1468,  -14'd1405,  14'd593,  -14'd581,  14'd2286,  -14'd1074,  -14'd169,  14'd1665,  14'd433,  -14'd1003,  -14'd1007,  14'd187,  
14'd767,  14'd1431,  -14'd1080,  -14'd4,  -14'd795,  14'd1499,  14'd324,  -14'd705,  -14'd1107,  -14'd456,  -14'd737,  14'd22,  14'd261,  14'd1825,  14'd200,  14'd763,  
14'd111,  14'd68,  14'd1040,  -14'd61,  14'd270,  -14'd1559,  -14'd211,  -14'd545,  14'd543,  -14'd197,  -14'd134,  14'd586,  14'd544,  14'd1723,  -14'd870,  14'd750,  
14'd261,  14'd1622,  -14'd1689,  -14'd514,  14'd215,  -14'd235,  14'd1073,  -14'd496,  14'd1017,  14'd1008,  14'd772,  14'd1120,  -14'd405,  14'd1699,  14'd309,  14'd28,  
-14'd778,  -14'd568,  14'd1327,  -14'd171,  14'd317,  14'd92,  14'd1016,  14'd1352,  -14'd349,  14'd1260,  14'd1084,  -14'd261,  14'd578,  14'd630,  -14'd337,  14'd137,  
-14'd1055,  -14'd543,  14'd1008,  -14'd352,  -14'd1161,  14'd275,  14'd767,  14'd303,  -14'd114,  14'd780,  14'd159,  -14'd223,  14'd623,  -14'd683,  14'd6,  -14'd1435,  
14'd143,  14'd1198,  -14'd79,  -14'd838,  14'd223,  -14'd870,  14'd593,  -14'd1174,  14'd146,  -14'd2,  -14'd752,  14'd1578,  14'd1410,  -14'd317,  14'd135,  -14'd220,  
14'd845,  14'd729,  -14'd802,  14'd443,  14'd275,  -14'd54,  14'd274,  -14'd2030,  14'd145,  -14'd2102,  -14'd966,  14'd556,  -14'd84,  14'd1059,  -14'd770,  14'd530,  
-14'd114,  14'd664,  -14'd2050,  -14'd760,  14'd1251,  -14'd704,  14'd810,  -14'd746,  14'd746,  -14'd343,  14'd814,  14'd799,  14'd1252,  -14'd593,  14'd95,  -14'd392,  
14'd508,  14'd46,  14'd367,  14'd1056,  -14'd1068,  -14'd240,  14'd1047,  14'd128,  -14'd32,  14'd832,  14'd725,  -14'd234,  14'd183,  14'd647,  14'd1442,  14'd993,  
14'd435,  14'd25,  14'd441,  -14'd417,  -14'd120,  -14'd156,  14'd1113,  14'd830,  14'd838,  14'd569,  14'd1384,  -14'd503,  14'd167,  -14'd1481,  14'd192,  -14'd442,  
14'd1396,  -14'd1516,  14'd863,  14'd1845,  14'd802,  14'd1027,  -14'd1591,  14'd457,  14'd121,  14'd964,  14'd231,  14'd1023,  14'd901,  14'd1401,  14'd1049,  14'd798,  
14'd1197,  -14'd1953,  -14'd1022,  -14'd760,  14'd1141,  -14'd389,  14'd665,  -14'd1069,  -14'd798,  -14'd382,  -14'd1033,  14'd658,  14'd1135,  14'd413,  -14'd251,  -14'd860,  
14'd343,  -14'd1276,  -14'd834,  14'd112,  -14'd596,  14'd5,  -14'd888,  -14'd1212,  14'd10,  14'd1057,  -14'd724,  14'd618,  -14'd487,  14'd1049,  -14'd177,  14'd1334,  
14'd472,  -14'd77,  14'd512,  -14'd710,  14'd1193,  -14'd1491,  14'd1708,  -14'd107,  -14'd781,  14'd55,  14'd123,  14'd594,  14'd615,  14'd41,  -14'd64,  14'd1151,  
14'd740,  -14'd1005,  -14'd1214,  -14'd4,  -14'd871,  14'd236,  14'd701,  14'd341,  14'd1427,  14'd1278,  -14'd897,  -14'd746,  -14'd505,  14'd1298,  -14'd202,  14'd471,  
-14'd692,  14'd927,  -14'd556,  14'd700,  -14'd775,  14'd508,  14'd350,  -14'd255,  -14'd62,  -14'd880,  14'd1175,  14'd989,  14'd395,  -14'd1101,  -14'd593,  14'd137,  
-14'd173,  -14'd903,  -14'd411,  14'd485,  14'd1703,  -14'd173,  -14'd103,  -14'd11,  -14'd248,  -14'd368,  14'd1119,  -14'd746,  -14'd232,  -14'd369,  -14'd162,  -14'd1061,  
-14'd343,  -14'd942,  -14'd941,  14'd644,  14'd1871,  14'd165,  14'd411,  14'd308,  14'd418,  14'd1309,  14'd29,  14'd1109,  14'd296,  -14'd783,  -14'd409,  14'd1225,  
14'd842,  14'd1564,  -14'd481,  -14'd1411,  -14'd236,  -14'd843,  -14'd27,  -14'd528,  -14'd1783,  -14'd1099,  14'd129,  -14'd60,  -14'd228,  14'd959,  14'd1,  -14'd1103,  
-14'd677,  -14'd627,  14'd1803,  14'd105,  -14'd433,  -14'd953,  -14'd1320,  14'd789,  -14'd1597,  -14'd1442,  -14'd1504,  -14'd588,  -14'd677,  14'd3077,  -14'd605,  -14'd395,  
-14'd611,  14'd749,  14'd450,  -14'd227,  14'd341,  14'd3,  -14'd1,  -14'd170,  -14'd706,  -14'd1030,  -14'd84,  -14'd444,  -14'd225,  14'd1252,  14'd1208,  -14'd1120,  
-14'd1079,  -14'd873,  -14'd1216,  -14'd919,  -14'd818,  14'd1469,  -14'd496,  14'd332,  -14'd518,  -14'd931,  14'd786,  14'd233,  14'd663,  14'd1709,  14'd2002,  14'd1608,  
-14'd2222,  14'd971,  14'd155,  14'd1344,  -14'd307,  -14'd427,  14'd83,  -14'd133,  -14'd1521,  -14'd215,  14'd1116,  14'd630,  -14'd691,  -14'd206,  14'd1976,  14'd631
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule



module bias_fc2_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC2-1][0:`OUTPUT_NUM_FC2-1][`WD_BIAS:0] weight	 = {
		24'd376858,  24'd432250,  24'd29999,  -24'd21180,  24'd203900,  -24'd35257,  24'd214653,  -24'd285062,  24'd149942,  24'd172424,  24'd241287,  24'd324760,  24'd306054,  24'd109385,  24'd386902,  24'd1789,  
24'd28800,  24'd347429,  24'd509845,  24'd403218,  24'd55283,  24'd293083,  -24'd21746,  -24'd254371,  -24'd400996,  -24'd132702,  -24'd107502,  -24'd140243,  -24'd206663,  -24'd140441,  24'd143746,  24'd39439,  
24'd236044,  24'd268803,  24'd150150,  24'd385287,  -24'd213047,  24'd26023,  -24'd343539,  24'd332436,  -24'd397889,  -24'd209506,  -24'd133163,  24'd243649,  -24'd9532,  24'd307082,  -24'd132963,  -24'd159572,  
-24'd53911,  24'd55608,  -24'd63297,  24'd287278,  24'd231376,  24'd227915,  -24'd149391,  24'd406123,  -24'd279679,  24'd37076,  24'd251134,  24'd110896,  -24'd132970,  24'd307661,  24'd327144,  24'd66815,  
24'd131364,  24'd119973,  -24'd302322,  24'd158931,  24'd47008,  -24'd154135,  -24'd42487,  24'd329397,  24'd366838,  24'd373655,  24'd391455,  24'd142308,  24'd61661,  24'd27682,  24'd173948,  -24'd11642,  
24'd233626,  -24'd79977,  24'd87200,  24'd305044
	 };
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule


module wieght_fc2_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2*`OUTPUT_BATCH_FC2)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC1*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC2*`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2-1][0:`OUTPUT_NUM_FC2-1][0:`OUTPUT_NUM_FC1-1][`WD:0] weight	 = {
14'd168,  -14'd674,  -14'd1094,  14'd1558,  14'd2074,  -14'd421,  14'd870,  14'd1633,  -14'd1381,  -14'd256,  -14'd1566,  14'd1621,  -14'd1118,  -14'd377,  14'd1870,  14'd582,  
14'd868,  -14'd119,  -14'd78,  14'd935,  14'd1023,  -14'd1907,  14'd125,  14'd1935,  14'd84,  -14'd196,  -14'd471,  -14'd185,  -14'd684,  14'd567,  14'd416,  -14'd858,  
14'd763,  14'd1327,  -14'd1039,  14'd597,  -14'd370,  14'd335,  14'd519,  14'd1427,  -14'd358,  -14'd1447,  14'd401,  14'd687,  14'd1196,  14'd325,  -14'd1720,  -14'd656,  
-14'd401,  14'd382,  14'd307,  14'd767,  -14'd754,  14'd537,  -14'd1231,  14'd97,  14'd993,  -14'd1026,  14'd64,  -14'd602,  14'd136,  14'd1379,  -14'd346,  14'd929,  
14'd105,  14'd1083,  14'd676,  -14'd798,  -14'd244,  -14'd902,  -14'd443,  14'd225,  14'd696,  14'd1764,  -14'd872,  -14'd1169,  14'd745,  -14'd368,  -14'd1072,  14'd894,  
-14'd253,  -14'd156,  14'd445,  14'd67,  14'd634,  -14'd1342,  -14'd991,  14'd258,  -14'd1173,  14'd546,  -14'd1395,  -14'd1285,  14'd754,  14'd517,  14'd1351,  -14'd661,  
-14'd97,  -14'd847,  -14'd297,  14'd2439,  -14'd323,  -14'd952,  14'd123,  -14'd254,  -14'd1163,  -14'd623,  -14'd1520,  14'd1706,  -14'd986,  -14'd953,  14'd439,  14'd869,  
14'd741,  14'd319,  -14'd1197,  -14'd58,  14'd769,  -14'd159,  -14'd1435,  -14'd943,  
-14'd723,  -14'd920,  14'd297,  14'd92,  -14'd145,  -14'd803,  -14'd1449,  -14'd1645,  14'd270,  14'd227,  14'd376,  -14'd1799,  14'd16,  14'd299,  14'd1365,  14'd831,  
-14'd54,  -14'd517,  14'd1357,  -14'd588,  -14'd107,  14'd1387,  14'd317,  -14'd667,  14'd303,  -14'd1242,  -14'd407,  -14'd680,  14'd728,  14'd865,  14'd818,  14'd41,  
-14'd426,  -14'd165,  14'd1692,  14'd725,  14'd407,  14'd270,  -14'd303,  -14'd97,  14'd1104,  -14'd1513,  14'd583,  14'd289,  14'd675,  -14'd41,  -14'd990,  -14'd1580,  
14'd370,  -14'd1439,  -14'd130,  14'd424,  14'd1591,  14'd900,  -14'd1386,  -14'd573,  -14'd632,  14'd945,  -14'd821,  14'd875,  14'd1346,  14'd572,  14'd314,  14'd274,  
14'd497,  14'd142,  14'd352,  14'd50,  -14'd886,  14'd164,  -14'd1011,  14'd68,  -14'd1356,  -14'd803,  14'd153,  -14'd259,  -14'd725,  -14'd1052,  14'd414,  -14'd535,  
14'd72,  -14'd144,  14'd1259,  -14'd374,  -14'd70,  -14'd997,  -14'd68,  14'd46,  -14'd31,  -14'd147,  -14'd1005,  14'd921,  14'd1182,  14'd868,  -14'd1134,  14'd412,  
14'd1306,  14'd1238,  -14'd756,  14'd181,  14'd755,  -14'd395,  14'd741,  -14'd2228,  14'd1092,  14'd177,  -14'd826,  -14'd1495,  -14'd118,  14'd701,  -14'd1389,  14'd1204,  
14'd214,  -14'd91,  -14'd677,  -14'd43,  14'd1005,  14'd290,  14'd1409,  -14'd449,  
-14'd1310,  -14'd646,  14'd657,  14'd949,  -14'd215,  14'd842,  14'd210,  14'd506,  -14'd940,  14'd28,  14'd75,  -14'd513,  14'd166,  14'd765,  -14'd71,  14'd767,  
-14'd962,  14'd393,  -14'd830,  14'd140,  14'd318,  14'd821,  -14'd258,  14'd479,  -14'd1129,  -14'd1076,  -14'd549,  14'd701,  -14'd234,  14'd436,  -14'd313,  14'd1286,  
-14'd519,  14'd1154,  14'd1001,  14'd1073,  -14'd1072,  14'd1374,  -14'd329,  14'd866,  14'd1430,  14'd575,  -14'd551,  -14'd466,  -14'd385,  14'd1607,  14'd299,  -14'd937,  
14'd133,  -14'd1415,  14'd1579,  14'd240,  14'd185,  -14'd1967,  14'd1218,  14'd525,  -14'd90,  14'd975,  14'd1133,  14'd1055,  14'd890,  -14'd483,  -14'd1223,  -14'd286,  
-14'd800,  14'd158,  -14'd173,  -14'd569,  -14'd41,  -14'd678,  -14'd198,  14'd837,  -14'd255,  14'd640,  14'd1046,  -14'd773,  -14'd1399,  -14'd627,  14'd389,  -14'd1167,  
14'd611,  -14'd1262,  -14'd1474,  -14'd371,  14'd886,  14'd397,  14'd1069,  14'd566,  14'd83,  -14'd851,  14'd391,  -14'd741,  -14'd1510,  14'd1721,  14'd635,  -14'd51,  
-14'd1148,  -14'd52,  14'd37,  -14'd81,  -14'd638,  14'd631,  -14'd1117,  14'd1194,  14'd114,  14'd890,  14'd496,  14'd372,  -14'd324,  -14'd51,  14'd1059,  14'd561,  
14'd197,  14'd87,  14'd123,  -14'd202,  14'd1922,  -14'd729,  -14'd62,  14'd677,  
14'd572,  -14'd149,  14'd367,  -14'd60,  14'd932,  14'd384,  14'd381,  -14'd991,  -14'd1422,  14'd72,  -14'd1480,  -14'd1043,  14'd654,  14'd254,  14'd337,  14'd509,  
14'd1317,  14'd608,  -14'd419,  -14'd1219,  14'd611,  14'd687,  14'd1140,  14'd185,  14'd790,  -14'd1308,  14'd53,  -14'd2150,  14'd438,  14'd15,  14'd1092,  14'd2062,  
14'd260,  14'd24,  14'd325,  14'd244,  14'd1452,  -14'd543,  -14'd1628,  14'd898,  -14'd576,  14'd387,  14'd703,  -14'd1716,  14'd1020,  14'd515,  -14'd2188,  -14'd604,  
-14'd391,  14'd1309,  14'd1467,  14'd126,  -14'd378,  14'd229,  14'd76,  -14'd49,  14'd831,  14'd1165,  -14'd41,  14'd36,  14'd463,  -14'd717,  14'd337,  -14'd1320,  
-14'd413,  14'd197,  -14'd431,  14'd1306,  -14'd1633,  14'd123,  -14'd1866,  -14'd35,  14'd813,  -14'd1409,  -14'd183,  14'd744,  -14'd1544,  -14'd555,  14'd1187,  14'd378,  
-14'd484,  -14'd726,  14'd813,  -14'd260,  -14'd1081,  14'd443,  14'd306,  -14'd973,  -14'd494,  -14'd392,  14'd1076,  -14'd667,  14'd517,  -14'd55,  14'd1272,  -14'd303,  
14'd1093,  -14'd120,  14'd279,  -14'd535,  14'd1320,  14'd1819,  -14'd263,  -14'd3420,  14'd233,  -14'd562,  -14'd737,  -14'd487,  14'd113,  -14'd2228,  -14'd1033,  14'd1411,  
14'd99,  14'd95,  14'd140,  -14'd1406,  -14'd1588,  -14'd700,  14'd278,  14'd1463,  
-14'd782,  -14'd150,  -14'd1056,  -14'd607,  14'd751,  14'd999,  14'd764,  -14'd378,  -14'd360,  14'd793,  -14'd1534,  14'd833,  14'd771,  14'd605,  14'd306,  14'd52,  
14'd576,  -14'd150,  14'd795,  -14'd828,  -14'd87,  14'd1032,  14'd594,  14'd83,  14'd513,  -14'd1230,  -14'd188,  14'd908,  14'd317,  -14'd514,  14'd737,  -14'd578,  
-14'd897,  14'd911,  -14'd481,  -14'd154,  -14'd138,  14'd39,  -14'd323,  14'd1646,  -14'd1643,  -14'd127,  -14'd2370,  -14'd545,  14'd436,  14'd801,  14'd1663,  14'd967,  
14'd891,  -14'd1230,  -14'd1332,  14'd1302,  14'd188,  14'd1194,  14'd491,  -14'd728,  -14'd378,  -14'd203,  14'd680,  -14'd405,  -14'd68,  14'd1054,  14'd648,  -14'd663,  
14'd1341,  -14'd546,  14'd745,  -14'd1399,  14'd1936,  -14'd338,  -14'd508,  14'd1205,  14'd43,  -14'd5,  -14'd790,  -14'd12,  14'd323,  14'd139,  -14'd450,  14'd1147,  
-14'd52,  -14'd766,  14'd1178,  -14'd1242,  -14'd411,  -14'd345,  -14'd299,  14'd155,  -14'd1271,  14'd659,  14'd505,  14'd490,  14'd872,  -14'd1050,  -14'd351,  -14'd252,  
-14'd467,  14'd276,  14'd634,  -14'd1682,  -14'd44,  14'd4,  14'd886,  -14'd705,  -14'd267,  -14'd62,  -14'd661,  14'd2770,  14'd756,  -14'd440,  -14'd1474,  -14'd293,  
14'd1541,  -14'd677,  14'd1234,  -14'd786,  -14'd396,  14'd869,  14'd69,  -14'd777,  
-14'd1444,  -14'd67,  14'd1332,  14'd105,  -14'd1608,  14'd1622,  14'd557,  -14'd1226,  -14'd290,  14'd815,  14'd2202,  -14'd1238,  -14'd776,  14'd9,  -14'd377,  -14'd150,  
-14'd154,  -14'd76,  -14'd738,  14'd594,  14'd338,  14'd897,  14'd1186,  -14'd29,  -14'd114,  14'd203,  14'd904,  -14'd43,  -14'd666,  14'd1164,  -14'd1005,  -14'd171,  
-14'd819,  14'd391,  14'd195,  -14'd348,  14'd874,  14'd427,  -14'd952,  -14'd1500,  14'd718,  14'd160,  -14'd474,  14'd1406,  -14'd1508,  14'd42,  -14'd297,  14'd449,  
14'd1052,  14'd263,  14'd751,  14'd1278,  14'd1597,  14'd264,  14'd1747,  14'd202,  -14'd2118,  14'd306,  -14'd800,  -14'd213,  14'd1280,  14'd201,  14'd925,  -14'd1188,  
-14'd430,  -14'd1201,  -14'd1091,  14'd530,  -14'd1518,  14'd969,  -14'd88,  -14'd109,  14'd275,  14'd1112,  14'd445,  14'd626,  -14'd1142,  14'd209,  -14'd388,  14'd621,  
14'd702,  -14'd381,  14'd308,  -14'd1657,  14'd590,  14'd1668,  14'd505,  -14'd856,  -14'd139,  14'd63,  14'd905,  14'd151,  -14'd118,  14'd658,  14'd364,  14'd842,  
14'd1013,  14'd575,  14'd987,  -14'd391,  14'd928,  -14'd955,  14'd1374,  14'd980,  14'd165,  -14'd670,  14'd193,  -14'd431,  -14'd991,  14'd15,  14'd1223,  -14'd519,  
-14'd46,  14'd1143,  14'd2181,  14'd1128,  -14'd424,  -14'd1138,  -14'd876,  -14'd318,  
14'd485,  -14'd701,  14'd797,  -14'd618,  -14'd1047,  -14'd1360,  -14'd1800,  14'd739,  -14'd1874,  -14'd527,  -14'd1333,  -14'd942,  -14'd671,  14'd831,  -14'd1221,  14'd553,  
-14'd359,  14'd269,  14'd43,  -14'd379,  14'd708,  -14'd1212,  -14'd187,  14'd740,  14'd826,  14'd910,  14'd819,  -14'd775,  -14'd269,  14'd189,  -14'd346,  14'd1293,  
-14'd482,  14'd667,  14'd1274,  14'd359,  14'd1897,  -14'd519,  -14'd1626,  -14'd1341,  14'd4,  -14'd708,  -14'd305,  -14'd122,  -14'd1276,  -14'd440,  -14'd1088,  -14'd3177,  
14'd332,  14'd297,  -14'd44,  14'd783,  14'd234,  14'd600,  14'd669,  14'd816,  14'd882,  14'd539,  14'd343,  14'd1322,  14'd1134,  -14'd2398,  -14'd456,  14'd278,  
14'd251,  14'd272,  -14'd1097,  -14'd815,  -14'd1682,  14'd1574,  -14'd203,  14'd241,  -14'd957,  14'd77,  14'd167,  -14'd760,  14'd817,  14'd825,  14'd553,  14'd221,  
-14'd481,  -14'd1374,  -14'd128,  14'd687,  -14'd631,  -14'd1203,  -14'd784,  -14'd366,  -14'd534,  14'd734,  14'd64,  -14'd812,  14'd535,  14'd1157,  -14'd1234,  14'd1672,  
-14'd581,  -14'd898,  -14'd468,  -14'd565,  -14'd570,  14'd190,  14'd1608,  14'd400,  -14'd1040,  -14'd1260,  -14'd40,  14'd657,  -14'd534,  -14'd712,  -14'd493,  14'd448,  
-14'd484,  14'd708,  -14'd1617,  -14'd396,  14'd1180,  14'd502,  14'd51,  -14'd442,  
14'd863,  -14'd255,  -14'd806,  -14'd950,  14'd957,  14'd526,  -14'd1141,  -14'd285,  -14'd497,  -14'd524,  -14'd1341,  14'd725,  14'd920,  -14'd182,  14'd1430,  14'd208,  
14'd491,  14'd567,  -14'd473,  14'd85,  -14'd1200,  14'd592,  -14'd477,  14'd1914,  14'd462,  14'd1668,  -14'd551,  -14'd1255,  14'd1469,  -14'd197,  14'd674,  14'd502,  
14'd620,  -14'd131,  -14'd392,  14'd188,  14'd1390,  -14'd266,  14'd1034,  -14'd103,  -14'd771,  -14'd577,  14'd112,  -14'd1182,  14'd1513,  14'd647,  -14'd277,  -14'd1343,  
14'd249,  14'd686,  14'd675,  -14'd1733,  -14'd180,  14'd483,  14'd1457,  14'd358,  14'd86,  14'd844,  -14'd931,  14'd722,  14'd582,  14'd750,  14'd429,  -14'd672,  
14'd27,  14'd860,  14'd967,  -14'd305,  14'd405,  -14'd1865,  14'd1504,  14'd352,  14'd2084,  -14'd1315,  -14'd170,  -14'd1908,  14'd446,  -14'd491,  14'd314,  14'd616,  
-14'd160,  -14'd1112,  -14'd1483,  14'd1166,  -14'd607,  -14'd148,  14'd256,  -14'd188,  -14'd1811,  -14'd1256,  14'd1374,  14'd246,  14'd1617,  -14'd1344,  -14'd149,  -14'd723,  
-14'd592,  14'd807,  -14'd700,  14'd1431,  14'd376,  -14'd856,  -14'd1172,  -14'd373,  -14'd799,  14'd500,  -14'd316,  14'd315,  -14'd979,  -14'd381,  -14'd142,  14'd1117,  
-14'd1046,  -14'd616,  -14'd46,  14'd871,  14'd553,  14'd1165,  -14'd58,  14'd835,  
14'd262,  14'd679,  -14'd911,  -14'd153,  -14'd1083,  14'd522,  -14'd1450,  -14'd95,  -14'd654,  -14'd967,  -14'd711,  14'd970,  -14'd309,  14'd1933,  -14'd186,  14'd201,  
14'd269,  -14'd1888,  14'd919,  14'd1210,  14'd437,  14'd1318,  14'd52,  -14'd786,  14'd63,  -14'd945,  -14'd665,  14'd71,  -14'd495,  14'd566,  -14'd1827,  -14'd308,  
-14'd162,  14'd691,  -14'd568,  -14'd394,  14'd94,  14'd760,  -14'd1528,  14'd412,  -14'd951,  14'd560,  -14'd867,  -14'd626,  14'd628,  14'd1094,  -14'd708,  14'd399,  
14'd331,  14'd729,  -14'd374,  14'd231,  14'd1188,  14'd632,  -14'd1052,  14'd107,  -14'd673,  14'd874,  14'd1397,  14'd317,  -14'd1563,  14'd817,  14'd1459,  14'd1354,  
14'd781,  -14'd843,  14'd389,  -14'd877,  14'd804,  14'd278,  14'd176,  -14'd1062,  14'd1060,  14'd1134,  -14'd598,  14'd205,  -14'd660,  -14'd681,  14'd356,  -14'd427,  
14'd656,  -14'd1015,  14'd489,  -14'd106,  -14'd1011,  -14'd209,  -14'd645,  14'd191,  -14'd437,  -14'd643,  -14'd121,  14'd285,  14'd563,  -14'd268,  -14'd599,  -14'd1078,  
14'd159,  -14'd302,  14'd1990,  -14'd857,  14'd338,  -14'd1553,  -14'd148,  -14'd430,  14'd936,  -14'd614,  -14'd1583,  14'd315,  -14'd540,  -14'd206,  -14'd267,  14'd914,  
14'd977,  14'd674,  14'd921,  14'd502,  -14'd1369,  -14'd573,  14'd645,  14'd1646,  
-14'd1012,  14'd149,  -14'd487,  14'd243,  14'd777,  14'd178,  14'd704,  14'd2377,  -14'd780,  14'd412,  14'd976,  -14'd259,  -14'd361,  -14'd603,  14'd650,  -14'd353,  
-14'd311,  14'd1007,  14'd786,  -14'd829,  14'd274,  -14'd570,  14'd768,  -14'd319,  14'd474,  14'd741,  -14'd163,  14'd470,  14'd151,  14'd1306,  14'd573,  -14'd592,  
-14'd586,  14'd1649,  -14'd869,  14'd543,  -14'd52,  -14'd2580,  -14'd911,  14'd1232,  -14'd1932,  -14'd653,  14'd495,  14'd1672,  14'd2776,  14'd1226,  -14'd128,  -14'd512,  
14'd1242,  14'd384,  14'd1363,  -14'd1180,  14'd84,  -14'd816,  -14'd3795,  -14'd652,  14'd948,  14'd642,  -14'd223,  14'd2041,  14'd175,  -14'd456,  -14'd489,  14'd2150,  
14'd581,  -14'd235,  -14'd666,  -14'd747,  -14'd1277,  14'd405,  -14'd491,  14'd756,  -14'd926,  -14'd232,  14'd996,  -14'd395,  14'd840,  -14'd247,  -14'd103,  -14'd619,  
-14'd1213,  14'd1906,  14'd139,  -14'd541,  -14'd299,  14'd1189,  -14'd420,  -14'd456,  -14'd953,  14'd689,  -14'd169,  14'd101,  14'd1046,  -14'd191,  14'd37,  14'd210,  
14'd277,  -14'd210,  -14'd1083,  -14'd348,  14'd196,  -14'd2559,  14'd94,  -14'd1317,  14'd311,  -14'd684,  -14'd323,  14'd105,  14'd583,  -14'd5,  -14'd858,  14'd1666,  
-14'd1087,  14'd1240,  -14'd917,  14'd207,  14'd1447,  14'd674,  -14'd200,  14'd680,  
-14'd792,  14'd1636,  -14'd916,  14'd574,  14'd1074,  14'd1063,  -14'd662,  -14'd438,  -14'd336,  14'd370,  -14'd3826,  -14'd474,  14'd1152,  14'd239,  14'd1354,  14'd1869,  
-14'd53,  -14'd322,  -14'd2438,  -14'd1235,  14'd527,  14'd336,  14'd746,  14'd1286,  14'd640,  -14'd1623,  -14'd1837,  -14'd1374,  14'd1066,  14'd173,  14'd2086,  14'd580,  
14'd344,  14'd1168,  14'd1505,  14'd1244,  -14'd1227,  14'd500,  14'd242,  14'd262,  -14'd63,  -14'd837,  14'd1428,  -14'd407,  -14'd592,  14'd371,  14'd632,  -14'd2239,  
-14'd353,  -14'd1200,  -14'd1146,  14'd130,  -14'd108,  14'd1442,  -14'd1207,  14'd1550,  14'd877,  14'd1358,  -14'd2511,  14'd1196,  -14'd532,  14'd977,  14'd622,  14'd6,  
14'd596,  -14'd379,  14'd1162,  14'd217,  14'd17,  -14'd980,  14'd12,  14'd1161,  -14'd528,  -14'd403,  -14'd824,  -14'd685,  14'd296,  14'd1249,  -14'd1440,  -14'd643,  
14'd683,  -14'd93,  14'd963,  -14'd115,  -14'd2489,  -14'd137,  -14'd553,  14'd730,  -14'd1225,  -14'd591,  14'd113,  14'd928,  14'd1489,  -14'd1112,  -14'd1462,  -14'd183,  
-14'd77,  -14'd1243,  -14'd886,  -14'd292,  -14'd791,  14'd2171,  -14'd25,  -14'd1420,  -14'd808,  14'd1408,  14'd1280,  14'd1352,  14'd635,  -14'd1653,  -14'd720,  14'd232,  
-14'd1012,  -14'd615,  14'd420,  -14'd886,  -14'd319,  -14'd95,  14'd687,  14'd1209,  
14'd270,  14'd574,  -14'd1256,  14'd236,  14'd1619,  14'd1444,  -14'd334,  -14'd253,  -14'd98,  14'd1920,  14'd642,  14'd1064,  -14'd21,  14'd390,  -14'd250,  14'd2113,  
14'd1223,  -14'd610,  -14'd301,  -14'd372,  -14'd127,  -14'd494,  14'd1547,  14'd1222,  14'd103,  14'd1902,  -14'd554,  14'd753,  -14'd646,  14'd951,  14'd920,  -14'd1358,  
-14'd891,  -14'd958,  14'd72,  14'd457,  -14'd144,  14'd1107,  14'd477,  14'd373,  -14'd1753,  14'd775,  -14'd205,  14'd736,  14'd1652,  14'd247,  -14'd736,  14'd86,  
-14'd223,  -14'd129,  -14'd718,  14'd1596,  14'd1541,  14'd2082,  14'd1262,  14'd1521,  -14'd1289,  -14'd826,  14'd57,  14'd982,  14'd1296,  -14'd243,  14'd735,  14'd174,  
14'd3058,  -14'd302,  -14'd358,  -14'd556,  14'd414,  -14'd726,  14'd1423,  14'd1057,  14'd2159,  14'd1107,  -14'd1540,  14'd491,  -14'd1072,  -14'd1821,  -14'd481,  14'd78,  
-14'd213,  -14'd1169,  -14'd1617,  -14'd182,  -14'd125,  14'd898,  14'd171,  14'd217,  -14'd794,  -14'd712,  14'd1497,  14'd303,  14'd578,  -14'd1855,  -14'd332,  14'd199,  
-14'd155,  -14'd641,  14'd921,  14'd1993,  -14'd1698,  14'd2411,  14'd347,  -14'd452,  14'd467,  14'd963,  14'd1286,  14'd622,  -14'd186,  14'd374,  14'd101,  14'd410,  
14'd1020,  -14'd200,  14'd248,  -14'd1390,  14'd493,  -14'd894,  -14'd650,  -14'd26,  
14'd448,  14'd200,  14'd154,  -14'd130,  14'd584,  14'd731,  -14'd198,  -14'd1185,  -14'd835,  14'd434,  -14'd1671,  14'd37,  14'd1161,  14'd490,  -14'd588,  14'd490,  
14'd788,  14'd1609,  -14'd885,  -14'd422,  14'd96,  -14'd734,  14'd1329,  -14'd789,  -14'd265,  -14'd2202,  14'd18,  -14'd20,  14'd1221,  14'd427,  -14'd465,  -14'd144,  
-14'd744,  14'd432,  14'd1635,  -14'd525,  -14'd2085,  14'd1611,  -14'd288,  -14'd1403,  14'd526,  -14'd993,  -14'd1673,  14'd633,  -14'd498,  14'd73,  14'd1391,  14'd1132,  
-14'd119,  -14'd2535,  14'd1266,  -14'd596,  14'd396,  -14'd1722,  -14'd80,  -14'd622,  14'd1653,  -14'd116,  14'd1076,  -14'd85,  -14'd617,  -14'd1152,  -14'd936,  -14'd423,  
14'd1392,  14'd539,  14'd1166,  14'd1676,  -14'd785,  -14'd858,  -14'd1519,  14'd794,  -14'd1158,  14'd1312,  14'd726,  14'd1136,  14'd1125,  14'd1406,  -14'd447,  14'd295,  
14'd72,  -14'd575,  -14'd945,  -14'd360,  14'd1132,  14'd1037,  14'd1206,  14'd241,  14'd586,  -14'd85,  14'd1316,  14'd918,  -14'd170,  14'd24,  14'd1615,  14'd1702,  
-14'd842,  14'd302,  14'd703,  14'd960,  -14'd611,  14'd958,  14'd446,  14'd1083,  14'd579,  14'd467,  14'd1378,  -14'd359,  -14'd496,  -14'd684,  14'd1055,  -14'd849,  
14'd215,  -14'd799,  14'd718,  14'd1320,  14'd431,  -14'd184,  -14'd1262,  14'd109,  
14'd2517,  -14'd579,  14'd268,  14'd284,  14'd2097,  -14'd1094,  -14'd1882,  -14'd2151,  -14'd21,  -14'd202,  -14'd639,  -14'd1168,  14'd642,  14'd674,  14'd386,  14'd891,  
14'd2311,  14'd1389,  -14'd398,  -14'd171,  -14'd826,  14'd906,  14'd1044,  14'd2281,  14'd658,  -14'd351,  -14'd817,  -14'd1645,  -14'd967,  14'd695,  14'd51,  14'd19,  
14'd1771,  -14'd42,  -14'd625,  14'd1041,  14'd1618,  14'd2351,  14'd641,  -14'd1142,  14'd318,  14'd919,  -14'd72,  -14'd499,  -14'd386,  -14'd336,  14'd601,  -14'd2249,  
14'd16,  14'd576,  -14'd1200,  14'd690,  14'd1326,  -14'd225,  14'd854,  14'd1662,  14'd406,  -14'd113,  -14'd70,  14'd866,  14'd1113,  -14'd319,  -14'd969,  -14'd407,  
14'd911,  14'd522,  -14'd768,  14'd104,  -14'd752,  14'd721,  -14'd917,  -14'd1424,  14'd739,  -14'd1606,  14'd1066,  -14'd1746,  -14'd312,  14'd139,  -14'd649,  14'd1133,  
14'd1219,  -14'd8,  -14'd313,  14'd1486,  14'd144,  14'd11,  -14'd150,  14'd1682,  -14'd335,  14'd173,  14'd1240,  -14'd762,  -14'd705,  14'd603,  -14'd828,  14'd322,  
14'd797,  14'd405,  -14'd464,  -14'd1555,  -14'd877,  14'd753,  14'd990,  14'd1190,  -14'd812,  14'd475,  14'd1189,  -14'd1667,  14'd1195,  14'd1510,  -14'd699,  14'd1282,  
-14'd1377,  -14'd354,  -14'd776,  -14'd61,  -14'd176,  -14'd225,  14'd650,  14'd388,  
14'd196,  -14'd447,  14'd1162,  -14'd356,  14'd533,  -14'd400,  14'd699,  -14'd1712,  -14'd805,  14'd470,  -14'd1484,  -14'd1054,  14'd1186,  14'd155,  14'd2167,  -14'd282,  
14'd1160,  14'd797,  -14'd1468,  14'd335,  14'd83,  -14'd611,  14'd413,  14'd1558,  14'd621,  -14'd255,  14'd285,  -14'd1823,  14'd338,  -14'd1234,  14'd736,  14'd2179,  
14'd1028,  -14'd186,  14'd330,  14'd317,  14'd1125,  14'd941,  14'd845,  -14'd448,  14'd129,  -14'd937,  -14'd110,  -14'd369,  14'd1112,  -14'd1367,  -14'd1012,  -14'd1963,  
-14'd711,  -14'd1066,  -14'd891,  14'd2157,  -14'd328,  14'd1216,  -14'd1262,  14'd579,  14'd23,  14'd203,  -14'd1173,  14'd1477,  -14'd654,  -14'd729,  14'd750,  -14'd810,  
-14'd249,  14'd278,  14'd1514,  14'd1249,  -14'd346,  -14'd1114,  14'd860,  14'd258,  -14'd915,  -14'd609,  -14'd980,  14'd255,  14'd461,  -14'd1152,  14'd1155,  -14'd534,  
14'd13,  -14'd219,  -14'd865,  14'd833,  14'd23,  -14'd1258,  14'd1114,  14'd480,  -14'd967,  14'd760,  14'd673,  -14'd361,  14'd1265,  14'd183,  14'd389,  -14'd588,  
14'd560,  -14'd360,  -14'd1128,  -14'd435,  -14'd752,  14'd2217,  14'd680,  14'd31,  -14'd326,  14'd415,  14'd921,  -14'd24,  14'd199,  -14'd1198,  -14'd838,  14'd2351,  
14'd650,  -14'd536,  -14'd1511,  14'd1447,  14'd1715,  -14'd82,  14'd1054,  -14'd351,  
14'd65,  14'd363,  -14'd1092,  -14'd424,  -14'd109,  -14'd372,  -14'd120,  -14'd284,  14'd1543,  -14'd1737,  -14'd15,  -14'd88,  14'd797,  14'd925,  -14'd40,  14'd1166,  
14'd107,  -14'd284,  14'd1392,  14'd288,  -14'd1030,  -14'd204,  -14'd1598,  14'd468,  -14'd968,  -14'd1243,  -14'd326,  -14'd773,  -14'd695,  14'd584,  -14'd862,  -14'd445,  
14'd830,  14'd694,  14'd310,  -14'd524,  -14'd1342,  14'd1009,  -14'd973,  -14'd7,  -14'd506,  14'd1427,  14'd64,  14'd402,  14'd12,  -14'd394,  -14'd720,  14'd106,  
-14'd85,  14'd31,  14'd511,  -14'd401,  14'd898,  14'd382,  -14'd173,  14'd581,  -14'd511,  14'd85,  -14'd532,  14'd447,  -14'd967,  -14'd727,  -14'd340,  -14'd94,  
-14'd1282,  -14'd547,  14'd864,  14'd98,  -14'd1152,  -14'd830,  14'd957,  14'd785,  14'd279,  -14'd482,  -14'd585,  14'd937,  14'd6,  -14'd414,  -14'd1077,  14'd444,  
14'd1548,  14'd703,  -14'd24,  -14'd560,  14'd1066,  -14'd842,  14'd316,  14'd926,  14'd196,  14'd772,  14'd108,  -14'd571,  -14'd522,  -14'd84,  14'd758,  -14'd567,  
14'd956,  -14'd1308,  14'd596,  14'd217,  -14'd749,  14'd383,  -14'd749,  -14'd621,  -14'd508,  -14'd328,  -14'd427,  -14'd941,  -14'd985,  -14'd437,  14'd297,  14'd268,  
-14'd193,  14'd395,  14'd512,  14'd230,  14'd163,  -14'd460,  -14'd624,  -14'd1098,  
-14'd1119,  -14'd305,  14'd365,  -14'd337,  -14'd250,  14'd134,  14'd624,  14'd536,  14'd296,  -14'd244,  14'd417,  14'd633,  -14'd886,  -14'd576,  14'd969,  -14'd270,  
-14'd1072,  14'd947,  14'd607,  14'd782,  14'd459,  14'd439,  14'd329,  -14'd166,  -14'd648,  14'd544,  14'd182,  -14'd740,  -14'd1212,  14'd827,  14'd576,  14'd798,  
-14'd127,  14'd538,  14'd180,  -14'd157,  14'd1727,  -14'd399,  -14'd414,  -14'd551,  14'd1540,  -14'd1124,  14'd544,  14'd503,  14'd1085,  14'd813,  14'd742,  14'd1099,  
14'd316,  -14'd106,  14'd817,  -14'd664,  14'd212,  14'd1855,  -14'd915,  14'd794,  -14'd1288,  -14'd209,  -14'd396,  -14'd670,  14'd329,  14'd1559,  14'd564,  14'd662,  
-14'd118,  14'd24,  -14'd263,  14'd388,  14'd604,  14'd1187,  14'd1331,  14'd584,  14'd159,  -14'd1260,  14'd466,  -14'd135,  14'd119,  14'd490,  14'd98,  14'd1273,  
14'd1090,  14'd1293,  -14'd283,  14'd1583,  14'd790,  -14'd799,  14'd39,  -14'd1507,  -14'd355,  -14'd1161,  -14'd664,  14'd216,  14'd1251,  -14'd973,  14'd116,  -14'd512,  
14'd1577,  14'd615,  -14'd820,  -14'd778,  -14'd846,  -14'd1571,  14'd362,  -14'd38,  -14'd610,  -14'd730,  -14'd566,  -14'd1460,  -14'd276,  14'd440,  -14'd1365,  14'd381,  
14'd92,  -14'd146,  14'd513,  14'd502,  -14'd1018,  14'd137,  14'd5,  14'd1077,  
-14'd1137,  14'd721,  14'd73,  -14'd82,  14'd1670,  -14'd646,  -14'd145,  -14'd2634,  14'd572,  14'd461,  14'd278,  -14'd329,  -14'd425,  -14'd857,  -14'd1367,  -14'd1333,  
14'd64,  14'd781,  -14'd343,  14'd1307,  14'd220,  14'd961,  -14'd1549,  14'd939,  14'd427,  14'd321,  14'd1960,  14'd335,  14'd610,  14'd317,  14'd605,  -14'd1382,  
-14'd467,  -14'd412,  -14'd189,  -14'd811,  -14'd1309,  14'd801,  14'd983,  -14'd837,  14'd1514,  -14'd210,  -14'd155,  14'd736,  -14'd144,  14'd408,  14'd1593,  14'd804,  
14'd56,  14'd120,  -14'd1132,  -14'd101,  14'd1914,  14'd1232,  -14'd1986,  14'd398,  -14'd28,  14'd685,  14'd490,  -14'd953,  -14'd20,  14'd1336,  14'd94,  -14'd367,  
-14'd377,  -14'd227,  -14'd301,  -14'd697,  14'd460,  14'd557,  14'd189,  -14'd937,  14'd123,  -14'd551,  -14'd259,  14'd245,  14'd1552,  -14'd889,  -14'd328,  -14'd89,  
-14'd147,  14'd1492,  14'd57,  14'd1560,  -14'd973,  -14'd558,  -14'd889,  -14'd219,  14'd507,  14'd899,  14'd1113,  -14'd672,  -14'd1037,  14'd458,  14'd144,  -14'd900,  
14'd594,  -14'd610,  -14'd1478,  14'd551,  -14'd291,  -14'd719,  14'd252,  -14'd2978,  -14'd610,  14'd1027,  14'd965,  14'd1445,  14'd1047,  -14'd2115,  14'd254,  14'd304,  
14'd432,  -14'd278,  -14'd668,  -14'd783,  14'd204,  -14'd790,  -14'd680,  -14'd1168,  
-14'd803,  -14'd73,  14'd1318,  -14'd1262,  14'd332,  -14'd451,  14'd256,  -14'd827,  14'd403,  14'd1218,  14'd1007,  -14'd467,  -14'd114,  -14'd34,  14'd654,  14'd1100,  
-14'd495,  14'd99,  14'd1565,  14'd204,  -14'd380,  14'd1138,  14'd237,  -14'd1723,  -14'd1014,  14'd291,  -14'd755,  -14'd770,  14'd1102,  -14'd329,  14'd657,  -14'd1221,  
14'd584,  -14'd797,  14'd1238,  14'd1347,  -14'd1604,  -14'd265,  -14'd335,  14'd1610,  -14'd1361,  -14'd1296,  -14'd458,  14'd1464,  14'd1286,  14'd630,  14'd1168,  14'd83,  
-14'd312,  14'd433,  -14'd1654,  -14'd1481,  -14'd748,  14'd1389,  -14'd2508,  14'd344,  14'd1456,  14'd132,  -14'd305,  14'd622,  -14'd636,  14'd94,  -14'd587,  14'd658,  
14'd338,  14'd1324,  -14'd614,  14'd93,  14'd570,  14'd763,  14'd113,  -14'd25,  14'd434,  14'd877,  14'd569,  14'd1784,  14'd600,  14'd370,  14'd212,  14'd776,  
14'd301,  -14'd885,  -14'd948,  14'd69,  -14'd750,  -14'd970,  14'd530,  14'd20,  14'd846,  -14'd607,  -14'd344,  -14'd799,  -14'd990,  14'd775,  -14'd402,  -14'd519,  
14'd1154,  14'd682,  -14'd650,  14'd1763,  14'd496,  -14'd2,  14'd264,  -14'd816,  -14'd283,  14'd927,  -14'd766,  -14'd767,  14'd1270,  -14'd1864,  14'd932,  -14'd231,  
14'd1588,  -14'd145,  14'd593,  14'd75,  14'd269,  -14'd1028,  -14'd1445,  -14'd54,  
-14'd2080,  -14'd132,  -14'd1429,  -14'd250,  -14'd615,  14'd671,  14'd629,  -14'd1278,  14'd490,  14'd356,  14'd1348,  -14'd777,  14'd776,  -14'd778,  14'd529,  -14'd804,  
-14'd923,  -14'd117,  -14'd36,  14'd1707,  -14'd704,  -14'd635,  14'd784,  -14'd2012,  -14'd565,  14'd96,  14'd44,  14'd2055,  14'd726,  -14'd1440,  14'd1455,  -14'd80,  
14'd262,  -14'd620,  14'd287,  14'd80,  -14'd800,  -14'd7,  -14'd637,  14'd580,  14'd1140,  14'd425,  -14'd1214,  14'd1583,  -14'd1558,  14'd8,  14'd1773,  -14'd640,  
14'd379,  14'd205,  14'd461,  14'd175,  -14'd119,  14'd219,  -14'd39,  -14'd715,  14'd1486,  -14'd1468,  14'd1388,  -14'd1749,  14'd767,  14'd1256,  14'd465,  -14'd615,  
14'd133,  14'd528,  -14'd308,  -14'd130,  14'd375,  -14'd873,  14'd1283,  14'd392,  -14'd12,  14'd881,  -14'd1272,  14'd1916,  -14'd1077,  14'd1741,  -14'd829,  14'd244,  
-14'd614,  14'd57,  14'd968,  14'd741,  -14'd81,  14'd1112,  -14'd496,  14'd281,  -14'd91,  14'd852,  -14'd774,  14'd981,  -14'd1159,  14'd790,  14'd798,  14'd237,  
-14'd713,  14'd1360,  -14'd1255,  14'd244,  14'd1031,  -14'd532,  -14'd338,  -14'd464,  14'd1291,  14'd25,  -14'd231,  14'd358,  -14'd383,  14'd1525,  14'd716,  14'd413,  
-14'd14,  -14'd278,  -14'd563,  14'd1772,  14'd240,  -14'd1528,  14'd1336,  -14'd1529,  
-14'd614,  -14'd1588,  14'd1021,  14'd348,  -14'd1556,  -14'd405,  -14'd23,  14'd1816,  -14'd1508,  -14'd1113,  -14'd670,  -14'd501,  -14'd1271,  -14'd103,  14'd78,  14'd662,  
-14'd342,  -14'd607,  -14'd934,  -14'd142,  -14'd742,  14'd405,  14'd703,  14'd239,  -14'd537,  14'd757,  14'd1067,  14'd170,  -14'd1085,  -14'd386,  -14'd1305,  14'd810,  
14'd281,  14'd1436,  -14'd332,  -14'd312,  14'd560,  -14'd185,  -14'd924,  -14'd390,  -14'd208,  14'd298,  14'd1298,  -14'd1086,  -14'd818,  -14'd939,  14'd616,  -14'd689,  
14'd896,  14'd662,  14'd418,  14'd85,  -14'd2131,  -14'd985,  14'd431,  -14'd1007,  -14'd1080,  14'd1556,  14'd36,  -14'd782,  -14'd794,  14'd270,  14'd2772,  -14'd464,  
-14'd276,  -14'd1974,  -14'd314,  -14'd1110,  -14'd424,  -14'd50,  14'd1474,  -14'd446,  -14'd529,  14'd323,  -14'd672,  -14'd116,  -14'd514,  14'd1137,  14'd26,  14'd861,  
14'd51,  -14'd1122,  14'd1413,  14'd1367,  -14'd665,  14'd896,  -14'd1097,  -14'd1287,  14'd1315,  -14'd430,  -14'd229,  -14'd635,  -14'd612,  14'd130,  14'd829,  14'd434,  
14'd224,  14'd437,  -14'd73,  -14'd132,  14'd1452,  14'd2023,  14'd488,  -14'd799,  14'd454,  14'd2206,  14'd880,  -14'd272,  -14'd483,  14'd3040,  -14'd1206,  14'd216,  
14'd510,  -14'd1718,  14'd1087,  -14'd275,  -14'd1232,  -14'd1283,  -14'd571,  -14'd755,  
14'd485,  -14'd639,  14'd1173,  14'd1450,  -14'd459,  -14'd460,  -14'd710,  -14'd299,  -14'd166,  14'd1656,  14'd449,  14'd228,  -14'd490,  14'd1804,  14'd1075,  14'd1657,  
-14'd407,  14'd743,  14'd382,  -14'd1340,  14'd1402,  14'd510,  -14'd596,  14'd319,  -14'd1413,  14'd243,  14'd373,  14'd540,  -14'd1029,  14'd714,  14'd371,  14'd1423,  
-14'd441,  14'd162,  14'd367,  -14'd414,  14'd384,  -14'd2328,  -14'd1154,  14'd143,  -14'd1827,  14'd920,  -14'd808,  -14'd810,  14'd1790,  14'd871,  14'd595,  -14'd1631,  
14'd560,  -14'd136,  -14'd102,  14'd134,  14'd450,  -14'd154,  -14'd982,  -14'd1625,  -14'd788,  14'd966,  14'd461,  14'd1782,  14'd856,  14'd179,  14'd737,  14'd1093,  
14'd702,  14'd754,  14'd614,  -14'd1594,  14'd848,  -14'd147,  14'd1638,  14'd756,  -14'd499,  -14'd1122,  -14'd1303,  -14'd408,  14'd1586,  -14'd716,  -14'd1019,  14'd403,  
14'd1179,  -14'd395,  14'd353,  14'd795,  14'd1053,  14'd1039,  -14'd847,  -14'd603,  -14'd221,  -14'd136,  -14'd427,  -14'd485,  -14'd1164,  14'd432,  14'd542,  -14'd139,  
14'd1098,  -14'd1855,  -14'd585,  -14'd599,  -14'd96,  -14'd1244,  14'd880,  -14'd2124,  -14'd93,  -14'd1654,  -14'd540,  -14'd543,  14'd593,  -14'd148,  -14'd289,  14'd896,  
14'd358,  -14'd1037,  -14'd833,  14'd791,  -14'd590,  -14'd1618,  14'd641,  14'd189,  
14'd106,  14'd401,  -14'd966,  14'd941,  -14'd605,  14'd1366,  14'd152,  -14'd825,  -14'd660,  -14'd1511,  -14'd1110,  -14'd1032,  14'd544,  -14'd362,  -14'd1115,  14'd803,  
-14'd313,  14'd366,  -14'd1373,  14'd330,  -14'd910,  14'd164,  14'd1007,  14'd316,  -14'd228,  14'd724,  -14'd1011,  -14'd1192,  -14'd347,  -14'd806,  -14'd1025,  -14'd8,  
-14'd542,  14'd44,  14'd636,  -14'd935,  -14'd292,  14'd707,  -14'd883,  -14'd874,  14'd679,  -14'd51,  -14'd301,  14'd73,  -14'd610,  14'd258,  -14'd1652,  -14'd52,  
14'd834,  -14'd1464,  -14'd118,  -14'd1081,  -14'd842,  -14'd244,  -14'd455,  -14'd74,  -14'd577,  14'd72,  -14'd1211,  14'd135,  -14'd807,  -14'd306,  14'd1597,  -14'd564,  
-14'd1479,  -14'd1315,  -14'd1433,  -14'd287,  -14'd677,  -14'd359,  14'd1019,  -14'd800,  -14'd754,  14'd311,  -14'd1006,  14'd1333,  -14'd565,  14'd150,  -14'd1163,  14'd323,  
-14'd648,  14'd1512,  -14'd221,  -14'd6,  -14'd659,  14'd182,  14'd446,  -14'd372,  14'd478,  -14'd1259,  14'd1014,  14'd1149,  -14'd8,  14'd212,  14'd246,  14'd0,  
-14'd888,  -14'd1311,  -14'd96,  -14'd1206,  -14'd1736,  -14'd68,  -14'd49,  14'd148,  -14'd1595,  -14'd678,  -14'd1349,  14'd512,  -14'd993,  -14'd293,  14'd198,  -14'd1334,  
-14'd1574,  14'd1010,  -14'd1040,  -14'd1341,  -14'd118,  -14'd80,  14'd1058,  14'd292,  
14'd942,  -14'd406,  -14'd1410,  14'd551,  14'd620,  -14'd744,  14'd82,  14'd261,  -14'd569,  14'd562,  14'd1204,  -14'd85,  14'd355,  -14'd751,  14'd390,  14'd37,  
-14'd1537,  14'd376,  14'd220,  -14'd770,  -14'd275,  -14'd704,  -14'd1034,  14'd471,  -14'd227,  -14'd462,  -14'd913,  14'd542,  -14'd403,  -14'd267,  -14'd399,  14'd367,  
14'd12,  -14'd1018,  14'd18,  14'd874,  -14'd1121,  -14'd296,  14'd185,  -14'd198,  -14'd246,  -14'd526,  -14'd871,  -14'd739,  14'd205,  -14'd366,  -14'd1163,  -14'd806,  
-14'd264,  -14'd245,  -14'd816,  -14'd50,  -14'd357,  -14'd588,  14'd711,  14'd234,  14'd109,  -14'd362,  -14'd644,  14'd1021,  14'd77,  -14'd863,  14'd850,  -14'd313,  
14'd918,  -14'd1879,  14'd129,  -14'd518,  14'd489,  -14'd657,  14'd367,  -14'd714,  -14'd289,  14'd932,  -14'd924,  14'd606,  -14'd75,  -14'd34,  -14'd551,  14'd687,  
-14'd295,  14'd792,  14'd805,  -14'd1528,  -14'd1232,  -14'd227,  -14'd919,  14'd818,  -14'd22,  -14'd1484,  14'd757,  -14'd588,  14'd576,  -14'd116,  14'd1188,  -14'd597,  
-14'd865,  -14'd953,  14'd106,  14'd714,  14'd279,  14'd231,  -14'd1771,  -14'd1052,  -14'd77,  -14'd1163,  -14'd514,  -14'd1395,  -14'd791,  -14'd338,  14'd235,  -14'd814,  
14'd165,  14'd50,  -14'd1318,  -14'd1278,  -14'd1244,  -14'd788,  -14'd830,  -14'd16,  
-14'd281,  14'd301,  -14'd864,  14'd3,  -14'd1036,  14'd1177,  14'd287,  14'd160,  -14'd150,  -14'd1634,  14'd1075,  -14'd252,  -14'd642,  14'd866,  -14'd864,  -14'd164,  
-14'd638,  -14'd806,  -14'd1796,  -14'd1017,  -14'd806,  -14'd1455,  -14'd173,  -14'd237,  -14'd303,  -14'd1180,  -14'd987,  -14'd1371,  -14'd461,  14'd777,  -14'd353,  -14'd1104,  
-14'd395,  -14'd1144,  14'd168,  -14'd113,  14'd1405,  -14'd1124,  -14'd100,  -14'd1272,  -14'd1387,  -14'd1666,  -14'd264,  -14'd592,  -14'd997,  14'd216,  -14'd685,  -14'd250,  
14'd908,  14'd201,  -14'd821,  -14'd1290,  14'd209,  14'd389,  -14'd1871,  14'd978,  14'd450,  14'd460,  -14'd554,  -14'd444,  -14'd110,  -14'd289,  -14'd127,  -14'd204,  
14'd1087,  -14'd1123,  -14'd222,  -14'd1362,  -14'd676,  -14'd124,  14'd757,  -14'd355,  -14'd436,  -14'd727,  -14'd832,  -14'd786,  -14'd591,  -14'd1321,  -14'd812,  -14'd1110,  
-14'd1019,  -14'd1141,  14'd44,  -14'd583,  14'd601,  -14'd784,  14'd161,  14'd181,  -14'd271,  14'd17,  -14'd296,  14'd307,  14'd311,  -14'd330,  14'd104,  -14'd164,  
-14'd2011,  -14'd1152,  14'd1155,  -14'd1703,  -14'd884,  -14'd456,  -14'd743,  14'd1072,  14'd242,  14'd245,  -14'd147,  -14'd878,  14'd273,  -14'd1146,  -14'd1055,  -14'd696,  
14'd266,  14'd225,  14'd196,  14'd114,  -14'd207,  14'd397,  14'd284,  -14'd275,  
14'd442,  -14'd567,  -14'd1246,  14'd367,  14'd111,  14'd1563,  -14'd84,  -14'd266,  -14'd110,  -14'd1086,  -14'd2,  14'd115,  -14'd1320,  -14'd1329,  14'd1206,  -14'd624,  
14'd362,  14'd1003,  14'd323,  -14'd399,  14'd946,  14'd540,  -14'd939,  -14'd301,  -14'd512,  14'd580,  14'd827,  -14'd594,  -14'd605,  -14'd494,  -14'd569,  14'd463,  
-14'd139,  14'd177,  -14'd840,  -14'd1218,  14'd435,  -14'd125,  14'd939,  -14'd350,  -14'd125,  -14'd1365,  -14'd528,  -14'd775,  -14'd450,  -14'd161,  -14'd1104,  -14'd363,  
14'd746,  14'd82,  -14'd983,  14'd1200,  14'd1230,  14'd411,  14'd1526,  -14'd659,  14'd194,  14'd144,  -14'd718,  -14'd102,  14'd518,  -14'd113,  14'd456,  14'd26,  
-14'd981,  -14'd1513,  14'd309,  -14'd1460,  -14'd164,  -14'd697,  -14'd280,  -14'd1244,  14'd952,  -14'd363,  14'd1133,  -14'd852,  14'd910,  14'd953,  -14'd431,  -14'd83,  
14'd494,  14'd1184,  14'd61,  -14'd14,  14'd155,  -14'd1575,  14'd307,  -14'd676,  14'd394,  14'd585,  -14'd1652,  -14'd637,  -14'd180,  -14'd53,  -14'd848,  -14'd434,  
-14'd392,  -14'd686,  -14'd1260,  14'd495,  -14'd265,  -14'd582,  -14'd1513,  -14'd312,  -14'd1331,  14'd718,  -14'd570,  -14'd543,  -14'd635,  -14'd177,  -14'd1069,  -14'd791,  
-14'd613,  -14'd710,  14'd845,  -14'd562,  14'd208,  -14'd164,  -14'd275,  -14'd1171,  
-14'd754,  -14'd630,  14'd466,  14'd502,  -14'd1955,  14'd1089,  14'd552,  -14'd67,  14'd745,  -14'd223,  -14'd889,  14'd745,  -14'd39,  14'd1152,  14'd1489,  -14'd443,  
-14'd2741,  -14'd591,  14'd1615,  -14'd1127,  14'd79,  -14'd1299,  14'd823,  14'd35,  14'd605,  -14'd279,  14'd2217,  -14'd842,  -14'd2525,  14'd550,  -14'd241,  -14'd292,  
-14'd806,  14'd1140,  -14'd2352,  -14'd733,  14'd331,  14'd2006,  14'd1751,  -14'd213,  14'd819,  -14'd642,  -14'd673,  -14'd814,  -14'd27,  14'd90,  -14'd209,  14'd734,  
-14'd883,  14'd832,  14'd950,  14'd193,  14'd199,  14'd90,  14'd301,  -14'd358,  14'd993,  14'd1212,  14'd88,  -14'd251,  -14'd2418,  -14'd1,  14'd1778,  -14'd565,  
14'd249,  -14'd1495,  14'd987,  14'd563,  14'd1389,  -14'd1090,  14'd3404,  -14'd78,  -14'd1717,  14'd275,  -14'd76,  14'd156,  -14'd268,  -14'd781,  -14'd1756,  -14'd1349,  
14'd573,  14'd669,  14'd234,  -14'd29,  14'd987,  -14'd1115,  -14'd819,  -14'd643,  14'd225,  14'd1903,  14'd529,  14'd177,  14'd148,  14'd463,  -14'd1370,  14'd516,  
14'd991,  -14'd727,  14'd2123,  14'd1513,  14'd862,  -14'd607,  -14'd1384,  14'd1339,  14'd827,  14'd1910,  -14'd1063,  -14'd2024,  -14'd734,  14'd94,  -14'd121,  -14'd294,  
14'd908,  14'd627,  14'd1571,  14'd1431,  -14'd1285,  14'd1081,  14'd1389,  14'd959,  
-14'd1338,  -14'd1106,  14'd937,  14'd375,  -14'd986,  -14'd1665,  -14'd944,  -14'd419,  14'd466,  14'd384,  -14'd455,  14'd853,  14'd61,  -14'd1532,  14'd607,  14'd39,  
-14'd349,  -14'd862,  -14'd1368,  -14'd1217,  -14'd890,  -14'd265,  -14'd467,  -14'd824,  14'd500,  -14'd82,  -14'd600,  14'd134,  -14'd250,  14'd328,  14'd1379,  14'd1021,  
14'd453,  -14'd600,  -14'd733,  14'd323,  -14'd136,  14'd438,  14'd108,  -14'd301,  -14'd146,  14'd399,  -14'd1828,  14'd574,  14'd343,  14'd702,  -14'd214,  -14'd124,  
-14'd601,  14'd772,  -14'd142,  -14'd722,  -14'd617,  14'd708,  -14'd150,  -14'd854,  -14'd1146,  14'd101,  -14'd567,  -14'd943,  -14'd236,  -14'd450,  -14'd210,  14'd819,  
-14'd25,  -14'd1398,  14'd506,  -14'd162,  -14'd893,  14'd277,  -14'd686,  -14'd102,  14'd627,  -14'd927,  -14'd212,  -14'd397,  14'd231,  14'd48,  -14'd97,  14'd156,  
-14'd148,  -14'd499,  -14'd438,  -14'd1022,  -14'd108,  14'd680,  14'd53,  -14'd1711,  14'd853,  14'd145,  -14'd162,  14'd562,  -14'd841,  -14'd1034,  14'd264,  -14'd321,  
14'd722,  14'd124,  -14'd674,  -14'd390,  -14'd1177,  -14'd147,  -14'd699,  14'd291,  -14'd86,  -14'd36,  -14'd730,  -14'd1803,  -14'd425,  14'd340,  14'd147,  14'd90,  
-14'd72,  14'd363,  -14'd526,  -14'd256,  -14'd559,  14'd1160,  -14'd529,  14'd374,  
14'd2348,  14'd173,  14'd453,  -14'd54,  -14'd491,  14'd392,  14'd408,  -14'd1356,  14'd1175,  -14'd5,  14'd493,  -14'd1766,  14'd25,  -14'd1180,  -14'd657,  14'd828,  
14'd643,  -14'd560,  14'd309,  14'd417,  14'd693,  14'd1220,  14'd174,  14'd1849,  14'd649,  14'd936,  14'd30,  14'd834,  -14'd723,  14'd1205,  14'd726,  14'd510,  
14'd495,  -14'd1016,  14'd847,  14'd1116,  14'd42,  14'd1313,  14'd1588,  -14'd1615,  -14'd592,  14'd1463,  -14'd1459,  -14'd884,  14'd319,  -14'd1267,  -14'd1579,  -14'd1405,  
-14'd315,  -14'd356,  14'd879,  -14'd1195,  14'd471,  14'd516,  14'd554,  -14'd247,  -14'd1247,  14'd678,  14'd790,  14'd413,  -14'd811,  -14'd123,  -14'd1020,  14'd15,  
14'd1405,  -14'd2089,  14'd1376,  14'd459,  -14'd139,  14'd1768,  -14'd559,  -14'd950,  -14'd913,  -14'd1396,  14'd55,  -14'd1733,  -14'd282,  -14'd584,  14'd1474,  -14'd380,  
-14'd411,  14'd339,  14'd1176,  -14'd31,  -14'd1788,  -14'd1215,  14'd601,  -14'd908,  -14'd429,  14'd916,  14'd991,  14'd738,  14'd1489,  14'd681,  14'd1025,  14'd1210,  
14'd1020,  14'd1815,  -14'd1393,  -14'd49,  -14'd160,  -14'd1083,  14'd763,  14'd2887,  14'd147,  -14'd1054,  14'd145,  -14'd1064,  14'd91,  14'd1982,  -14'd1104,  14'd339,  
14'd231,  -14'd1470,  -14'd985,  -14'd1391,  14'd1031,  -14'd884,  -14'd658,  -14'd239,  
-14'd1464,  -14'd657,  -14'd1017,  14'd219,  14'd72,  14'd505,  14'd5,  -14'd56,  -14'd751,  -14'd430,  14'd694,  14'd107,  -14'd813,  14'd946,  -14'd470,  14'd230,  
-14'd863,  -14'd418,  -14'd686,  -14'd13,  14'd1103,  -14'd72,  -14'd368,  -14'd258,  14'd256,  14'd241,  14'd977,  14'd983,  14'd641,  -14'd856,  -14'd240,  -14'd2274,  
-14'd270,  14'd109,  14'd902,  -14'd674,  14'd625,  14'd377,  -14'd1331,  14'd316,  -14'd520,  14'd1231,  -14'd160,  14'd66,  -14'd1908,  14'd971,  -14'd522,  14'd360,  
14'd854,  -14'd394,  14'd225,  14'd229,  -14'd863,  14'd1542,  14'd1865,  -14'd213,  14'd467,  -14'd444,  14'd1299,  -14'd1436,  14'd140,  14'd1444,  14'd1717,  -14'd1003,  
-14'd1048,  -14'd60,  14'd270,  -14'd47,  14'd697,  -14'd881,  -14'd414,  -14'd100,  14'd768,  -14'd600,  -14'd1234,  14'd278,  -14'd1457,  -14'd453,  -14'd1115,  14'd524,  
-14'd554,  14'd329,  14'd32,  -14'd1060,  14'd354,  14'd869,  14'd347,  -14'd74,  -14'd17,  14'd910,  14'd434,  14'd1613,  -14'd1655,  -14'd479,  14'd154,  14'd1069,  
-14'd470,  14'd569,  -14'd224,  14'd638,  14'd375,  14'd187,  -14'd968,  14'd98,  14'd142,  -14'd52,  -14'd58,  14'd173,  -14'd69,  14'd66,  14'd410,  -14'd1880,  
14'd996,  -14'd192,  14'd1105,  -14'd458,  14'd1401,  14'd869,  14'd449,  14'd391,  
14'd366,  14'd265,  -14'd1142,  -14'd172,  14'd2361,  -14'd38,  14'd488,  14'd2180,  -14'd131,  -14'd417,  14'd741,  14'd1189,  -14'd750,  -14'd1410,  -14'd475,  -14'd973,  
14'd2097,  14'd1024,  -14'd967,  14'd432,  14'd360,  -14'd50,  -14'd166,  14'd183,  14'd81,  14'd1415,  -14'd623,  14'd12,  -14'd940,  14'd1096,  14'd648,  -14'd1275,  
14'd426,  -14'd510,  -14'd628,  14'd231,  -14'd4,  -14'd456,  14'd276,  14'd666,  -14'd515,  -14'd730,  14'd1832,  -14'd545,  -14'd305,  14'd1268,  -14'd798,  14'd559,  
-14'd231,  14'd1304,  14'd421,  14'd1338,  14'd661,  14'd80,  -14'd750,  -14'd340,  -14'd894,  -14'd401,  -14'd639,  14'd880,  -14'd160,  14'd167,  -14'd243,  14'd640,  
14'd767,  14'd1116,  -14'd706,  14'd658,  14'd860,  14'd1016,  -14'd761,  14'd346,  14'd713,  14'd378,  14'd777,  -14'd448,  -14'd307,  14'd801,  -14'd929,  14'd454,  
-14'd1332,  14'd646,  -14'd727,  14'd2220,  14'd1053,  -14'd1051,  -14'd1001,  -14'd864,  -14'd457,  14'd1121,  -14'd1655,  -14'd464,  14'd668,  14'd1350,  -14'd141,  -14'd782,  
14'd440,  -14'd665,  -14'd934,  14'd1197,  14'd183,  -14'd1139,  -14'd855,  14'd1069,  14'd923,  -14'd758,  -14'd1262,  14'd1349,  -14'd279,  -14'd2134,  -14'd21,  -14'd849,  
-14'd504,  14'd1980,  -14'd1024,  14'd1052,  -14'd422,  14'd196,  -14'd198,  -14'd676,  
14'd1355,  14'd17,  -14'd698,  14'd343,  -14'd195,  14'd717,  -14'd1035,  14'd1494,  -14'd553,  -14'd275,  -14'd368,  -14'd1183,  -14'd688,  -14'd738,  -14'd1296,  14'd1416,  
14'd360,  -14'd1225,  -14'd291,  -14'd488,  14'd1315,  14'd495,  -14'd847,  -14'd599,  -14'd933,  14'd628,  -14'd1159,  -14'd476,  -14'd1520,  -14'd826,  14'd692,  -14'd717,  
-14'd49,  14'd206,  -14'd1,  -14'd1,  14'd551,  14'd512,  -14'd519,  14'd269,  14'd230,  14'd116,  -14'd1042,  14'd301,  -14'd440,  14'd694,  -14'd177,  14'd64,  
-14'd853,  -14'd331,  14'd133,  -14'd479,  -14'd1071,  -14'd823,  -14'd1158,  -14'd733,  -14'd500,  14'd29,  14'd688,  -14'd660,  14'd603,  14'd1217,  -14'd501,  -14'd53,  
-14'd533,  14'd978,  14'd340,  14'd818,  -14'd890,  -14'd108,  14'd849,  -14'd292,  14'd65,  14'd749,  -14'd266,  14'd1030,  -14'd212,  14'd424,  -14'd834,  14'd701,  
-14'd1250,  -14'd193,  -14'd271,  14'd479,  14'd506,  -14'd743,  -14'd1156,  14'd477,  -14'd228,  -14'd596,  -14'd606,  -14'd626,  -14'd37,  -14'd1036,  14'd938,  -14'd340,  
14'd556,  14'd70,  -14'd405,  -14'd348,  -14'd1,  -14'd370,  14'd877,  14'd1360,  -14'd78,  -14'd1431,  -14'd647,  14'd419,  14'd762,  14'd429,  -14'd447,  -14'd432,  
14'd197,  14'd1143,  14'd1136,  14'd94,  14'd324,  14'd781,  -14'd218,  14'd1408,  
14'd2345,  14'd176,  -14'd47,  14'd1111,  14'd1331,  14'd42,  -14'd234,  14'd681,  -14'd1453,  -14'd564,  -14'd107,  -14'd1088,  14'd13,  -14'd212,  14'd660,  14'd482,  
14'd509,  14'd827,  -14'd1572,  14'd896,  -14'd1329,  14'd74,  14'd521,  14'd1759,  -14'd1161,  14'd1496,  14'd469,  14'd1361,  -14'd1162,  14'd587,  -14'd93,  -14'd827,  
-14'd173,  -14'd708,  14'd209,  -14'd282,  14'd847,  14'd1014,  14'd1743,  -14'd48,  14'd1365,  -14'd206,  -14'd1211,  -14'd1635,  -14'd1052,  -14'd203,  -14'd1370,  14'd491,  
-14'd252,  14'd143,  -14'd1168,  -14'd945,  14'd1384,  14'd461,  -14'd385,  -14'd999,  14'd1615,  14'd1758,  -14'd142,  -14'd353,  14'd795,  14'd25,  -14'd1701,  14'd4,  
14'd119,  14'd1356,  14'd1338,  14'd749,  14'd1000,  14'd537,  14'd71,  -14'd245,  -14'd487,  14'd1925,  -14'd710,  -14'd544,  14'd1540,  14'd1250,  -14'd193,  14'd324,  
-14'd1211,  14'd1098,  -14'd306,  14'd107,  -14'd481,  14'd762,  -14'd560,  -14'd31,  -14'd38,  14'd1382,  -14'd194,  14'd1035,  14'd1815,  -14'd352,  14'd629,  -14'd440,  
14'd210,  -14'd143,  -14'd493,  14'd606,  -14'd1096,  14'd357,  14'd1446,  14'd1385,  -14'd1549,  -14'd34,  14'd331,  14'd342,  14'd517,  -14'd468,  14'd1489,  14'd890,  
-14'd1250,  14'd544,  14'd374,  -14'd322,  -14'd479,  14'd184,  14'd162,  14'd1831,  
-14'd2243,  -14'd756,  14'd1133,  14'd73,  -14'd631,  -14'd1054,  14'd587,  14'd2177,  14'd220,  14'd245,  -14'd716,  14'd2239,  -14'd30,  14'd817,  14'd1755,  -14'd1031,  
-14'd308,  14'd1077,  14'd396,  -14'd1370,  14'd410,  -14'd1672,  14'd18,  -14'd320,  -14'd467,  -14'd988,  14'd1726,  -14'd192,  -14'd29,  14'd1471,  -14'd359,  -14'd275,  
-14'd1152,  -14'd567,  -14'd386,  14'd351,  -14'd409,  -14'd1169,  14'd174,  14'd702,  14'd105,  -14'd957,  14'd1453,  14'd451,  14'd418,  14'd310,  14'd200,  14'd2018,  
-14'd1459,  14'd1000,  14'd1948,  -14'd2747,  -14'd807,  -14'd2209,  -14'd1220,  14'd716,  -14'd769,  -14'd484,  14'd947,  14'd146,  -14'd805,  14'd31,  14'd79,  14'd585,  
-14'd2465,  14'd934,  14'd655,  -14'd1424,  14'd393,  -14'd2532,  -14'd283,  14'd313,  -14'd96,  -14'd1173,  -14'd75,  -14'd459,  14'd2253,  -14'd254,  -14'd1013,  -14'd196,  
14'd104,  14'd1323,  -14'd302,  -14'd1067,  -14'd219,  14'd715,  14'd180,  14'd398,  -14'd477,  14'd699,  -14'd669,  14'd1282,  14'd233,  -14'd129,  14'd213,  14'd362,  
14'd910,  14'd48,  -14'd222,  -14'd474,  -14'd316,  -14'd2409,  -14'd169,  -14'd828,  14'd129,  -14'd1470,  -14'd1592,  -14'd32,  14'd778,  14'd200,  14'd994,  -14'd396,  
14'd807,  14'd709,  -14'd108,  14'd546,  -14'd43,  14'd174,  -14'd1413,  14'd1871,  
14'd560,  14'd10,  14'd1432,  -14'd629,  -14'd833,  14'd167,  14'd1161,  -14'd926,  14'd1902,  14'd785,  14'd333,  14'd451,  -14'd113,  -14'd1543,  -14'd958,  14'd1735,  
14'd882,  14'd15,  14'd1464,  14'd826,  -14'd429,  14'd1026,  14'd229,  14'd1043,  14'd853,  14'd792,  -14'd74,  -14'd469,  -14'd1219,  -14'd456,  -14'd1938,  -14'd1916,  
14'd1216,  -14'd620,  -14'd227,  -14'd173,  -14'd1182,  14'd1676,  14'd1908,  -14'd1168,  14'd893,  -14'd86,  14'd223,  14'd661,  -14'd1070,  -14'd97,  14'd117,  -14'd499,  
14'd403,  -14'd1544,  14'd65,  -14'd1241,  14'd259,  -14'd263,  14'd134,  14'd421,  -14'd1857,  14'd102,  14'd169,  -14'd614,  -14'd589,  -14'd484,  -14'd1578,  -14'd571,  
14'd2434,  -14'd1442,  -14'd422,  14'd920,  14'd1863,  14'd819,  -14'd1270,  14'd1273,  -14'd57,  -14'd234,  14'd1056,  14'd987,  -14'd1495,  -14'd527,  14'd181,  14'd784,  
-14'd1022,  14'd6,  -14'd753,  14'd281,  -14'd687,  14'd423,  -14'd700,  14'd1831,  14'd570,  14'd662,  -14'd730,  14'd435,  14'd788,  14'd269,  14'd539,  -14'd500,  
-14'd416,  -14'd531,  -14'd756,  -14'd69,  -14'd1326,  -14'd204,  14'd296,  14'd1358,  -14'd600,  14'd451,  14'd209,  -14'd1435,  14'd1094,  14'd355,  14'd500,  -14'd431,  
-14'd1214,  -14'd535,  -14'd938,  14'd90,  14'd757,  14'd533,  14'd44,  14'd919,  
14'd538,  -14'd55,  -14'd1784,  14'd348,  -14'd1391,  14'd394,  14'd272,  14'd686,  -14'd1408,  -14'd427,  -14'd392,  14'd81,  -14'd547,  14'd509,  14'd459,  14'd1787,  
14'd705,  -14'd677,  14'd1025,  -14'd840,  -14'd957,  -14'd950,  -14'd472,  -14'd957,  14'd494,  -14'd1500,  14'd275,  14'd300,  -14'd38,  14'd598,  -14'd244,  -14'd1506,  
-14'd1353,  14'd37,  -14'd1387,  14'd586,  14'd956,  -14'd734,  -14'd1063,  14'd473,  -14'd1349,  -14'd1819,  14'd39,  -14'd160,  14'd811,  -14'd141,  -14'd189,  14'd1012,  
14'd966,  -14'd2222,  14'd391,  -14'd891,  -14'd695,  -14'd1072,  14'd319,  14'd543,  -14'd1065,  14'd406,  -14'd43,  14'd564,  -14'd57,  -14'd1660,  -14'd1632,  -14'd121,  
14'd1095,  -14'd474,  14'd705,  14'd60,  -14'd1133,  14'd172,  14'd797,  -14'd313,  14'd33,  14'd1732,  -14'd1418,  -14'd1209,  14'd716,  -14'd473,  -14'd1483,  -14'd52,  
-14'd331,  -14'd991,  14'd1117,  -14'd1068,  -14'd1308,  14'd747,  14'd47,  14'd1227,  -14'd1673,  -14'd233,  -14'd781,  -14'd601,  14'd908,  -14'd248,  -14'd189,  14'd1168,  
14'd452,  -14'd1341,  14'd1310,  -14'd1170,  -14'd248,  -14'd2472,  -14'd917,  14'd279,  -14'd250,  -14'd796,  -14'd810,  -14'd523,  14'd326,  14'd748,  -14'd1077,  14'd1567,  
14'd1144,  -14'd451,  14'd782,  -14'd690,  14'd494,  14'd11,  14'd1199,  14'd1831,  
-14'd949,  -14'd381,  -14'd1069,  14'd140,  -14'd780,  -14'd1082,  14'd316,  14'd45,  14'd640,  -14'd1077,  -14'd778,  14'd629,  14'd163,  -14'd160,  14'd903,  -14'd718,  
-14'd294,  -14'd133,  14'd106,  14'd607,  14'd1092,  14'd407,  -14'd49,  14'd74,  -14'd215,  -14'd643,  -14'd70,  -14'd1193,  14'd479,  -14'd1520,  -14'd708,  -14'd541,  
14'd1118,  -14'd1734,  -14'd1777,  14'd900,  -14'd619,  -14'd1611,  -14'd102,  -14'd1245,  -14'd269,  14'd907,  -14'd669,  -14'd1054,  -14'd904,  14'd41,  -14'd1066,  14'd27,  
14'd649,  14'd620,  -14'd733,  -14'd313,  -14'd393,  14'd270,  14'd144,  -14'd503,  14'd811,  14'd264,  14'd221,  -14'd635,  -14'd1175,  14'd61,  -14'd251,  14'd1148,  
14'd287,  14'd13,  -14'd602,  -14'd186,  -14'd177,  -14'd6,  -14'd116,  14'd232,  14'd47,  -14'd480,  -14'd935,  14'd581,  -14'd673,  -14'd921,  -14'd748,  14'd869,  
14'd986,  -14'd904,  -14'd845,  14'd1583,  -14'd1023,  14'd575,  -14'd933,  -14'd811,  14'd837,  -14'd1227,  14'd332,  -14'd1648,  -14'd649,  -14'd9,  -14'd1440,  14'd73,  
14'd757,  -14'd973,  -14'd494,  14'd64,  -14'd518,  14'd867,  14'd558,  14'd424,  14'd785,  -14'd295,  14'd684,  14'd236,  14'd849,  -14'd1565,  -14'd135,  14'd214,  
-14'd578,  -14'd731,  -14'd391,  -14'd311,  -14'd1011,  -14'd364,  14'd907,  -14'd21,  
14'd201,  -14'd779,  -14'd1169,  14'd11,  -14'd233,  14'd332,  -14'd356,  -14'd1197,  14'd1040,  -14'd857,  14'd990,  -14'd816,  14'd655,  -14'd1398,  -14'd348,  14'd254,  
-14'd354,  14'd618,  -14'd100,  14'd216,  14'd531,  14'd773,  14'd950,  14'd327,  14'd1487,  14'd552,  14'd357,  -14'd378,  -14'd1563,  -14'd356,  14'd950,  14'd703,  
14'd1781,  14'd883,  14'd225,  -14'd273,  -14'd60,  14'd220,  14'd946,  -14'd814,  14'd929,  14'd1193,  -14'd548,  14'd1502,  -14'd302,  -14'd1172,  -14'd1506,  -14'd1930,  
-14'd182,  -14'd748,  -14'd445,  14'd1816,  14'd517,  14'd279,  14'd1390,  14'd719,  -14'd1083,  14'd1451,  14'd432,  14'd78,  14'd715,  14'd1008,  14'd134,  14'd68,  
14'd315,  -14'd1421,  14'd367,  14'd2945,  14'd373,  14'd170,  14'd429,  14'd1094,  14'd1517,  -14'd1121,  14'd249,  14'd266,  -14'd1802,  14'd557,  -14'd955,  -14'd1028,  
14'd1493,  14'd990,  -14'd487,  -14'd28,  14'd1222,  14'd74,  14'd1556,  -14'd45,  14'd558,  -14'd838,  14'd499,  -14'd353,  14'd883,  -14'd69,  -14'd553,  14'd1101,  
14'd987,  14'd1222,  -14'd1090,  -14'd333,  -14'd852,  14'd409,  -14'd287,  14'd1433,  -14'd1591,  14'd147,  14'd599,  -14'd2607,  14'd92,  14'd1666,  14'd85,  14'd534,  
-14'd556,  -14'd553,  -14'd442,  -14'd303,  14'd916,  -14'd265,  14'd1118,  14'd650,  
14'd837,  -14'd410,  14'd737,  -14'd442,  -14'd1406,  -14'd412,  14'd569,  14'd811,  14'd143,  -14'd121,  -14'd469,  -14'd515,  -14'd311,  -14'd586,  14'd334,  14'd1419,  
-14'd1006,  -14'd1131,  -14'd646,  -14'd957,  14'd87,  14'd570,  -14'd475,  -14'd283,  14'd16,  14'd195,  -14'd1439,  -14'd374,  14'd1649,  -14'd956,  -14'd139,  14'd1606,  
-14'd488,  14'd1061,  -14'd64,  14'd371,  -14'd434,  -14'd840,  -14'd1504,  14'd143,  14'd75,  14'd550,  14'd1815,  14'd357,  14'd0,  -14'd640,  14'd797,  -14'd612,  
14'd1068,  14'd1615,  14'd714,  -14'd74,  -14'd676,  -14'd1445,  14'd2119,  -14'd1490,  -14'd9,  14'd1257,  14'd761,  -14'd1507,  -14'd1100,  14'd404,  -14'd527,  -14'd5,  
14'd992,  14'd899,  14'd221,  14'd472,  -14'd21,  -14'd2231,  -14'd1078,  14'd843,  14'd1169,  -14'd2235,  14'd1474,  -14'd1886,  -14'd1938,  -14'd926,  -14'd157,  14'd193,  
-14'd119,  14'd941,  14'd361,  -14'd631,  14'd889,  14'd1276,  -14'd931,  -14'd325,  14'd464,  14'd243,  -14'd839,  14'd107,  14'd663,  14'd935,  -14'd1580,  14'd154,  
14'd478,  14'd1815,  -14'd690,  -14'd2229,  14'd1903,  -14'd1053,  -14'd1763,  -14'd811,  14'd1074,  -14'd743,  14'd267,  -14'd343,  14'd518,  14'd214,  14'd980,  -14'd19,  
-14'd753,  14'd957,  14'd1238,  14'd892,  14'd1051,  14'd1478,  14'd552,  -14'd971,  
-14'd1791,  14'd510,  -14'd405,  14'd395,  14'd49,  -14'd523,  14'd1135,  -14'd1632,  -14'd1898,  14'd0,  14'd705,  14'd1653,  14'd91,  14'd119,  -14'd45,  14'd465,  
-14'd1426,  14'd204,  14'd862,  -14'd162,  -14'd492,  -14'd377,  14'd835,  14'd31,  14'd791,  -14'd1834,  -14'd36,  14'd255,  14'd1109,  -14'd382,  14'd1152,  -14'd226,  
14'd321,  -14'd761,  14'd921,  14'd244,  -14'd1669,  14'd166,  14'd960,  14'd1306,  -14'd324,  -14'd696,  -14'd759,  -14'd1391,  14'd400,  14'd346,  14'd908,  -14'd316,  
-14'd266,  -14'd1453,  -14'd975,  14'd793,  -14'd694,  14'd198,  14'd869,  14'd475,  14'd652,  14'd93,  14'd1121,  14'd551,  -14'd140,  14'd978,  -14'd129,  -14'd785,  
14'd1312,  14'd1579,  14'd741,  14'd1565,  14'd253,  -14'd1401,  -14'd70,  14'd197,  14'd65,  -14'd793,  14'd343,  14'd1359,  14'd608,  14'd55,  14'd941,  14'd1257,  
14'd648,  14'd454,  14'd483,  -14'd1237,  -14'd1111,  14'd1268,  14'd1020,  14'd346,  -14'd559,  14'd1189,  14'd121,  14'd262,  -14'd1656,  -14'd900,  14'd291,  -14'd68,  
14'd127,  -14'd409,  14'd1792,  -14'd1080,  14'd330,  14'd549,  -14'd557,  -14'd1243,  -14'd223,  14'd1181,  14'd344,  -14'd779,  -14'd439,  14'd2069,  -14'd719,  -14'd898,  
14'd69,  -14'd1853,  14'd698,  14'd300,  14'd860,  14'd946,  14'd1749,  14'd1214,  
14'd345,  14'd214,  14'd716,  14'd230,  -14'd292,  14'd166,  14'd1118,  14'd346,  14'd215,  14'd196,  -14'd671,  14'd339,  14'd895,  14'd357,  -14'd752,  -14'd443,  
-14'd135,  -14'd1914,  -14'd157,  -14'd788,  -14'd1412,  14'd238,  14'd252,  14'd15,  -14'd307,  -14'd1201,  14'd164,  -14'd1510,  -14'd1078,  14'd459,  14'd1128,  -14'd233,  
14'd137,  -14'd1261,  -14'd1018,  -14'd370,  14'd1391,  -14'd1093,  -14'd1240,  -14'd25,  -14'd823,  14'd96,  14'd763,  -14'd822,  14'd995,  14'd252,  -14'd1543,  -14'd1288,  
14'd22,  -14'd1758,  -14'd1605,  14'd484,  14'd400,  -14'd631,  -14'd945,  14'd1184,  14'd134,  14'd1,  14'd141,  -14'd686,  -14'd841,  14'd46,  -14'd526,  -14'd1208,  
-14'd699,  -14'd195,  -14'd494,  14'd979,  -14'd1984,  -14'd398,  -14'd198,  -14'd963,  -14'd970,  -14'd42,  -14'd919,  14'd569,  14'd608,  14'd562,  14'd889,  14'd585,  
-14'd794,  14'd823,  -14'd917,  14'd494,  -14'd1705,  -14'd493,  -14'd985,  14'd494,  14'd367,  -14'd442,  -14'd765,  14'd299,  -14'd636,  -14'd441,  -14'd527,  -14'd1815,  
-14'd116,  -14'd822,  -14'd228,  -14'd797,  -14'd832,  14'd281,  -14'd1498,  -14'd1014,  14'd697,  -14'd584,  -14'd807,  14'd848,  14'd515,  14'd1110,  -14'd385,  14'd328,  
-14'd50,  14'd349,  14'd394,  14'd47,  14'd1164,  14'd617,  -14'd803,  14'd161,  
-14'd1323,  -14'd962,  -14'd32,  14'd319,  -14'd700,  -14'd543,  -14'd117,  -14'd427,  14'd1020,  -14'd817,  14'd1182,  14'd104,  -14'd367,  -14'd555,  14'd1029,  -14'd624,  
14'd292,  -14'd328,  -14'd1033,  -14'd1728,  -14'd500,  -14'd1521,  -14'd1016,  -14'd1799,  -14'd840,  -14'd728,  -14'd178,  -14'd669,  -14'd569,  -14'd1408,  -14'd179,  -14'd1044,  
-14'd152,  -14'd527,  -14'd53,  -14'd305,  -14'd854,  14'd65,  -14'd148,  -14'd345,  14'd760,  14'd666,  -14'd429,  14'd261,  -14'd921,  -14'd622,  -14'd1073,  -14'd225,  
-14'd601,  -14'd1555,  14'd45,  14'd24,  -14'd990,  -14'd801,  14'd934,  14'd1342,  -14'd171,  14'd1297,  14'd415,  -14'd1554,  -14'd1058,  -14'd939,  -14'd1235,  -14'd574,  
-14'd789,  -14'd1149,  14'd72,  14'd280,  14'd704,  14'd983,  -14'd134,  -14'd892,  -14'd1338,  14'd833,  14'd50,  14'd973,  14'd626,  14'd675,  -14'd1027,  -14'd1901,  
14'd486,  14'd727,  -14'd1317,  14'd614,  -14'd209,  14'd141,  -14'd99,  -14'd1639,  -14'd865,  14'd555,  14'd402,  -14'd330,  14'd349,  -14'd1660,  14'd634,  14'd566,  
14'd1298,  -14'd938,  14'd616,  -14'd817,  -14'd147,  -14'd1484,  -14'd734,  -14'd517,  -14'd1108,  14'd1278,  -14'd187,  -14'd1381,  -14'd1054,  14'd1073,  14'd145,  14'd494,  
-14'd557,  -14'd1918,  14'd751,  14'd744,  -14'd1377,  -14'd1208,  -14'd206,  -14'd591,  
-14'd1451,  -14'd190,  -14'd1482,  -14'd609,  -14'd1350,  -14'd247,  -14'd1009,  14'd360,  14'd975,  -14'd1054,  14'd386,  14'd138,  -14'd999,  -14'd39,  14'd87,  -14'd1740,  
-14'd201,  14'd729,  -14'd1742,  14'd380,  -14'd946,  14'd782,  14'd311,  -14'd45,  -14'd354,  14'd893,  14'd701,  14'd96,  14'd183,  14'd812,  14'd1652,  -14'd797,  
14'd1538,  -14'd154,  -14'd649,  -14'd703,  -14'd247,  -14'd446,  -14'd581,  14'd272,  14'd1062,  14'd208,  14'd1745,  14'd574,  14'd1097,  14'd589,  14'd955,  14'd439,  
-14'd204,  14'd338,  14'd1612,  14'd1131,  -14'd1691,  -14'd138,  14'd64,  -14'd1368,  14'd471,  14'd209,  -14'd337,  -14'd296,  -14'd1261,  14'd1003,  14'd611,  14'd265,  
-14'd1174,  14'd404,  -14'd764,  -14'd513,  14'd384,  -14'd961,  14'd42,  -14'd749,  14'd690,  -14'd2226,  -14'd274,  -14'd488,  -14'd1985,  14'd2029,  -14'd736,  14'd1597,  
-14'd268,  -14'd321,  14'd899,  -14'd502,  14'd898,  14'd1304,  -14'd479,  -14'd699,  -14'd280,  -14'd212,  14'd833,  14'd226,  -14'd352,  14'd831,  14'd137,  -14'd538,  
-14'd285,  14'd775,  -14'd924,  -14'd1921,  14'd1198,  -14'd1006,  -14'd1629,  14'd168,  14'd107,  14'd68,  14'd165,  -14'd1580,  14'd208,  14'd1273,  14'd444,  -14'd981,  
-14'd1071,  14'd611,  -14'd992,  -14'd404,  -14'd203,  14'd992,  -14'd151,  14'd109,  
-14'd62,  14'd716,  14'd1077,  -14'd1434,  -14'd581,  14'd320,  -14'd1100,  -14'd1439,  -14'd1085,  14'd1700,  -14'd558,  -14'd1419,  14'd1714,  14'd519,  14'd145,  -14'd786,  
-14'd50,  14'd1128,  -14'd490,  14'd1368,  14'd249,  14'd858,  -14'd110,  -14'd2583,  -14'd156,  14'd1127,  14'd793,  -14'd1554,  -14'd128,  -14'd940,  14'd91,  -14'd24,  
-14'd460,  14'd359,  14'd239,  14'd493,  -14'd938,  -14'd1310,  -14'd1282,  -14'd273,  14'd941,  -14'd317,  -14'd1378,  -14'd43,  -14'd461,  14'd84,  14'd124,  -14'd40,  
14'd813,  -14'd980,  14'd342,  -14'd1501,  14'd1861,  14'd234,  -14'd1989,  -14'd497,  14'd201,  14'd2230,  14'd713,  14'd80,  14'd1781,  -14'd468,  -14'd1197,  14'd485,  
-14'd1140,  -14'd83,  -14'd322,  14'd940,  14'd897,  -14'd1140,  -14'd509,  14'd1114,  -14'd1776,  -14'd1052,  14'd2011,  14'd1277,  14'd526,  -14'd1244,  14'd886,  14'd1333,  
14'd606,  -14'd965,  -14'd1035,  14'd28,  14'd314,  14'd1414,  14'd655,  -14'd576,  14'd485,  -14'd352,  -14'd919,  14'd443,  14'd525,  -14'd633,  -14'd1501,  14'd1270,  
14'd516,  -14'd134,  -14'd916,  -14'd1301,  14'd1823,  -14'd166,  14'd118,  14'd159,  -14'd929,  14'd1656,  14'd977,  -14'd1245,  -14'd532,  -14'd303,  -14'd642,  14'd603,  
14'd215,  -14'd925,  -14'd361,  -14'd487,  14'd1569,  -14'd481,  14'd1135,  14'd1787,  
14'd1115,  14'd306,  14'd1789,  -14'd405,  14'd718,  14'd500,  14'd1043,  -14'd1754,  14'd157,  -14'd270,  -14'd243,  -14'd984,  14'd1192,  -14'd263,  -14'd1566,  14'd1012,  
14'd367,  14'd1051,  -14'd1322,  -14'd718,  14'd580,  14'd23,  14'd1070,  14'd1603,  -14'd267,  14'd478,  -14'd535,  -14'd620,  -14'd464,  14'd622,  14'd344,  -14'd1488,  
-14'd299,  -14'd535,  -14'd1044,  -14'd1230,  14'd1584,  14'd644,  14'd876,  14'd559,  14'd428,  14'd453,  -14'd1128,  -14'd1273,  14'd487,  -14'd23,  14'd744,  14'd453,  
-14'd1081,  -14'd1437,  -14'd255,  -14'd527,  -14'd232,  14'd479,  14'd355,  14'd628,  -14'd2035,  14'd1332,  14'd470,  -14'd588,  14'd1251,  14'd518,  -14'd165,  14'd898,  
14'd1313,  -14'd1173,  14'd1877,  14'd325,  -14'd122,  -14'd1406,  14'd451,  -14'd515,  14'd989,  14'd493,  -14'd755,  -14'd1118,  -14'd1077,  -14'd65,  14'd353,  -14'd1441,  
14'd217,  14'd882,  -14'd1556,  -14'd245,  -14'd231,  -14'd98,  -14'd134,  14'd1118,  14'd667,  14'd2119,  14'd590,  -14'd381,  -14'd480,  14'd672,  -14'd1017,  -14'd4,  
-14'd53,  14'd266,  -14'd407,  -14'd173,  -14'd533,  14'd1163,  14'd978,  14'd1752,  -14'd666,  14'd1273,  14'd23,  -14'd562,  -14'd460,  14'd221,  14'd41,  -14'd265,  
-14'd860,  -14'd2255,  14'd1072,  14'd23,  14'd67,  -14'd138,  14'd75,  -14'd260,  
-14'd702,  14'd174,  14'd1960,  -14'd33,  -14'd1104,  -14'd194,  -14'd477,  -14'd787,  14'd137,  -14'd1130,  14'd729,  -14'd2129,  -14'd828,  -14'd99,  -14'd983,  14'd563,  
-14'd343,  14'd1801,  14'd1210,  14'd212,  -14'd825,  -14'd1122,  14'd187,  14'd2,  14'd1418,  14'd277,  14'd1667,  14'd199,  -14'd956,  14'd1256,  -14'd980,  -14'd1550,  
14'd1610,  14'd121,  14'd1152,  14'd1066,  -14'd1126,  -14'd267,  14'd232,  14'd581,  14'd767,  -14'd991,  -14'd1437,  14'd1062,  14'd1107,  -14'd621,  -14'd11,  -14'd278,  
14'd1315,  14'd27,  14'd478,  -14'd785,  -14'd608,  -14'd166,  -14'd992,  -14'd487,  -14'd1318,  -14'd328,  14'd266,  14'd900,  14'd628,  14'd209,  -14'd864,  14'd894,  
-14'd124,  -14'd804,  -14'd385,  -14'd996,  14'd1302,  14'd2214,  -14'd587,  14'd1504,  -14'd1187,  -14'd92,  14'd22,  -14'd442,  -14'd737,  -14'd710,  14'd293,  -14'd237,  
14'd956,  -14'd365,  -14'd595,  -14'd259,  14'd564,  -14'd347,  14'd834,  -14'd220,  14'd1276,  -14'd859,  14'd133,  -14'd776,  14'd1618,  14'd484,  14'd427,  14'd95,  
14'd662,  14'd321,  -14'd176,  14'd601,  -14'd579,  14'd263,  14'd151,  14'd1866,  14'd454,  -14'd923,  14'd714,  -14'd1208,  -14'd572,  14'd899,  14'd1045,  14'd1892,  
-14'd564,  -14'd431,  14'd1455,  14'd1309,  -14'd94,  -14'd682,  -14'd492,  14'd433,  
-14'd33,  14'd753,  14'd484,  -14'd573,  -14'd1148,  14'd703,  14'd460,  14'd373,  14'd120,  14'd69,  -14'd162,  -14'd313,  -14'd1003,  -14'd751,  -14'd203,  -14'd361,  
14'd647,  -14'd528,  14'd310,  -14'd496,  -14'd137,  -14'd1184,  14'd103,  -14'd445,  14'd110,  -14'd1261,  -14'd1644,  14'd28,  14'd396,  14'd220,  -14'd690,  -14'd887,  
-14'd954,  14'd1451,  14'd425,  -14'd729,  -14'd158,  -14'd1017,  -14'd575,  -14'd546,  14'd646,  -14'd252,  -14'd177,  -14'd120,  14'd725,  -14'd832,  -14'd545,  14'd376,  
14'd292,  -14'd772,  -14'd475,  14'd524,  14'd330,  -14'd351,  -14'd415,  -14'd906,  -14'd329,  14'd640,  14'd268,  -14'd559,  14'd1065,  -14'd1068,  -14'd244,  -14'd1275,  
-14'd889,  -14'd167,  14'd905,  14'd156,  14'd627,  -14'd93,  -14'd60,  -14'd90,  14'd504,  -14'd466,  14'd916,  14'd100,  -14'd249,  -14'd417,  -14'd325,  -14'd399,  
-14'd180,  -14'd273,  -14'd489,  14'd771,  14'd346,  -14'd1274,  -14'd340,  -14'd529,  -14'd709,  14'd901,  -14'd1340,  -14'd209,  -14'd612,  -14'd865,  14'd957,  -14'd58,  
14'd1058,  14'd51,  14'd170,  14'd161,  -14'd903,  -14'd1542,  -14'd143,  -14'd292,  -14'd1289,  -14'd307,  -14'd318,  -14'd1219,  -14'd331,  14'd90,  -14'd41,  14'd1153,  
-14'd760,  -14'd193,  14'd171,  -14'd310,  -14'd901,  14'd413,  14'd60,  -14'd1157,  
14'd33,  -14'd139,  -14'd303,  14'd958,  14'd221,  -14'd530,  -14'd1284,  14'd460,  -14'd1366,  -14'd650,  14'd4,  -14'd1209,  -14'd362,  -14'd582,  14'd123,  14'd14,  
-14'd229,  -14'd849,  -14'd763,  14'd274,  -14'd280,  -14'd78,  -14'd124,  -14'd1321,  -14'd76,  14'd518,  14'd807,  -14'd814,  14'd437,  -14'd839,  -14'd38,  14'd38,  
14'd363,  -14'd1697,  -14'd125,  -14'd1201,  -14'd1189,  14'd131,  14'd655,  -14'd273,  -14'd1059,  -14'd996,  14'd455,  -14'd37,  -14'd34,  -14'd582,  -14'd513,  -14'd74,  
14'd794,  14'd1022,  -14'd594,  14'd1238,  -14'd519,  -14'd1535,  -14'd307,  -14'd90,  -14'd1372,  14'd238,  14'd339,  -14'd1617,  -14'd171,  -14'd633,  14'd1401,  -14'd525,  
-14'd1470,  -14'd1143,  14'd607,  -14'd259,  -14'd515,  -14'd831,  14'd967,  -14'd696,  -14'd1092,  -14'd289,  -14'd600,  -14'd137,  -14'd359,  -14'd1630,  14'd347,  -14'd31,  
-14'd379,  -14'd185,  14'd561,  -14'd1027,  -14'd817,  14'd606,  -14'd675,  -14'd1367,  -14'd1352,  -14'd1362,  -14'd435,  -14'd595,  -14'd633,  14'd736,  14'd1533,  -14'd37,  
14'd558,  -14'd678,  -14'd1383,  -14'd102,  14'd1099,  14'd812,  14'd1070,  14'd430,  -14'd170,  14'd143,  -14'd186,  -14'd542,  14'd342,  14'd105,  -14'd1704,  -14'd833,  
-14'd1644,  -14'd1529,  14'd397,  -14'd1411,  -14'd674,  14'd311,  14'd298,  -14'd555,  
14'd37,  -14'd1399,  -14'd1180,  14'd771,  -14'd222,  14'd292,  -14'd249,  -14'd3204,  -14'd1489,  -14'd716,  -14'd464,  14'd1175,  -14'd162,  14'd407,  14'd852,  -14'd402,  
-14'd417,  -14'd257,  -14'd639,  -14'd294,  14'd283,  14'd435,  14'd967,  -14'd1216,  -14'd595,  14'd1863,  14'd1535,  14'd1236,  -14'd373,  14'd868,  14'd855,  14'd1125,  
14'd516,  14'd1766,  14'd1068,  14'd626,  14'd673,  -14'd475,  14'd919,  -14'd827,  14'd918,  14'd1449,  14'd107,  -14'd1278,  -14'd1741,  14'd764,  -14'd583,  -14'd1730,  
14'd820,  -14'd833,  14'd296,  -14'd1282,  14'd1268,  14'd1124,  14'd130,  -14'd43,  -14'd792,  14'd218,  14'd676,  14'd475,  14'd795,  -14'd226,  14'd813,  -14'd1303,  
14'd340,  14'd833,  -14'd561,  -14'd2163,  -14'd225,  -14'd186,  14'd1931,  -14'd649,  -14'd197,  -14'd864,  -14'd337,  -14'd1100,  14'd414,  -14'd63,  -14'd952,  -14'd552,  
14'd1162,  14'd344,  -14'd1085,  -14'd1233,  14'd1060,  -14'd739,  -14'd1416,  -14'd1060,  -14'd588,  14'd2122,  14'd242,  14'd1242,  14'd415,  -14'd714,  -14'd1073,  14'd408,  
-14'd716,  -14'd588,  -14'd260,  -14'd218,  -14'd185,  -14'd1787,  -14'd515,  -14'd1146,  14'd524,  -14'd414,  14'd1546,  -14'd534,  14'd274,  14'd2990,  -14'd96,  14'd1056,  
-14'd705,  14'd543,  14'd2023,  -14'd155,  -14'd119,  14'd548,  14'd359,  14'd38,  
14'd991,  -14'd215,  14'd855,  14'd777,  -14'd240,  -14'd1380,  -14'd251,  14'd116,  -14'd494,  14'd1360,  14'd2238,  14'd902,  -14'd1498,  -14'd1214,  -14'd1306,  14'd207,  
-14'd693,  -14'd546,  14'd1004,  14'd14,  -14'd307,  -14'd948,  14'd1127,  14'd928,  -14'd1040,  14'd260,  14'd554,  14'd1309,  -14'd1626,  -14'd331,  14'd391,  14'd123,  
14'd122,  -14'd54,  14'd419,  14'd507,  14'd118,  14'd900,  14'd221,  14'd207,  -14'd212,  14'd393,  14'd717,  -14'd538,  -14'd1583,  14'd52,  -14'd2825,  -14'd681,  
-14'd701,  14'd973,  -14'd14,  14'd1693,  -14'd2108,  14'd447,  14'd1504,  14'd1006,  14'd1287,  -14'd1866,  -14'd1080,  -14'd1520,  14'd1211,  -14'd984,  14'd822,  14'd521,  
14'd465,  -14'd341,  14'd343,  14'd1444,  14'd311,  14'd683,  14'd1173,  14'd569,  14'd182,  -14'd1327,  -14'd1115,  -14'd426,  -14'd1612,  -14'd2355,  -14'd292,  -14'd345,  
14'd762,  14'd54,  -14'd608,  -14'd1430,  14'd1911,  14'd197,  14'd77,  -14'd343,  14'd665,  14'd84,  14'd1646,  14'd667,  14'd108,  -14'd17,  -14'd1256,  14'd123,  
14'd395,  -14'd357,  14'd1871,  14'd2423,  -14'd661,  14'd2663,  -14'd241,  -14'd509,  14'd489,  -14'd440,  14'd500,  14'd473,  14'd315,  -14'd2002,  14'd799,  14'd619,  
14'd171,  -14'd856,  14'd572,  -14'd975,  -14'd326,  -14'd711,  14'd884,  -14'd518,  
-14'd146,  14'd587,  14'd348,  -14'd507,  14'd738,  -14'd704,  -14'd2,  14'd1617,  14'd2416,  -14'd1205,  14'd668,  -14'd1040,  -14'd1284,  -14'd1641,  -14'd691,  -14'd201,  
14'd749,  -14'd316,  -14'd581,  14'd1519,  -14'd134,  14'd444,  -14'd399,  -14'd340,  14'd30,  14'd451,  -14'd748,  -14'd875,  -14'd1196,  14'd317,  14'd1859,  14'd616,  
14'd266,  -14'd1126,  -14'd623,  14'd608,  14'd2091,  14'd521,  14'd65,  14'd1383,  14'd176,  14'd53,  14'd875,  -14'd1242,  14'd539,  14'd560,  -14'd22,  14'd238,  
-14'd410,  14'd575,  14'd14,  -14'd486,  14'd792,  -14'd28,  14'd26,  14'd450,  14'd252,  -14'd1196,  -14'd1564,  -14'd594,  14'd940,  14'd359,  14'd744,  14'd380,  
-14'd941,  14'd576,  -14'd283,  -14'd20,  -14'd466,  14'd893,  -14'd269,  14'd212,  14'd1665,  -14'd1073,  -14'd1199,  -14'd1809,  -14'd111,  14'd1290,  14'd787,  14'd1530,  
14'd1093,  14'd773,  -14'd693,  14'd2009,  -14'd157,  14'd387,  -14'd92,  14'd1179,  14'd1316,  14'd294,  -14'd925,  14'd982,  14'd1513,  -14'd569,  -14'd270,  -14'd244,  
-14'd318,  14'd613,  -14'd3027,  -14'd1293,  14'd530,  -14'd988,  -14'd1977,  14'd2213,  14'd950,  -14'd990,  -14'd751,  -14'd929,  -14'd118,  -14'd1320,  14'd264,  -14'd329,  
-14'd744,  14'd2273,  14'd967,  -14'd554,  -14'd492,  -14'd1069,  14'd60,  14'd385,  
14'd128,  -14'd594,  -14'd1913,  14'd565,  14'd1120,  14'd434,  -14'd250,  -14'd1001,  -14'd204,  14'd1720,  -14'd2053,  14'd574,  14'd634,  14'd557,  14'd1273,  -14'd999,  
14'd1483,  14'd537,  14'd1022,  14'd1517,  14'd1456,  14'd1132,  14'd967,  14'd261,  14'd206,  -14'd1577,  -14'd471,  14'd11,  14'd888,  -14'd599,  14'd1526,  -14'd1249,  
-14'd1317,  -14'd1190,  14'd975,  14'd245,  -14'd1212,  -14'd401,  14'd258,  14'd601,  14'd1733,  -14'd1272,  -14'd470,  14'd398,  14'd422,  14'd1331,  14'd1286,  14'd1671,  
14'd247,  -14'd1263,  14'd999,  -14'd1066,  14'd156,  -14'd56,  -14'd1543,  14'd321,  14'd217,  14'd305,  -14'd3,  14'd611,  -14'd467,  14'd200,  -14'd1640,  14'd716,  
-14'd1045,  14'd432,  14'd344,  14'd469,  14'd904,  -14'd1182,  -14'd386,  -14'd1175,  -14'd1069,  14'd934,  -14'd1119,  14'd1695,  14'd2116,  14'd1271,  -14'd430,  -14'd107,  
-14'd557,  14'd183,  -14'd1068,  -14'd936,  -14'd874,  14'd782,  14'd605,  14'd813,  14'd432,  -14'd519,  -14'd488,  14'd650,  14'd1500,  14'd1557,  14'd100,  -14'd337,  
14'd1268,  -14'd1595,  14'd857,  -14'd1403,  -14'd13,  14'd379,  -14'd1219,  -14'd1428,  14'd304,  14'd112,  -14'd1523,  14'd1231,  -14'd430,  -14'd2218,  14'd645,  14'd1101,  
-14'd647,  14'd444,  -14'd670,  14'd1241,  14'd1161,  14'd105,  -14'd804,  -14'd863,  
-14'd1456,  -14'd417,  -14'd778,  -14'd54,  -14'd265,  -14'd683,  14'd1395,  -14'd1843,  14'd2252,  14'd691,  14'd937,  -14'd744,  -14'd319,  14'd1080,  -14'd463,  14'd942,  
14'd684,  -14'd771,  14'd1360,  14'd885,  14'd73,  14'd1292,  14'd1549,  -14'd1570,  -14'd1338,  -14'd506,  -14'd856,  -14'd1015,  14'd1677,  -14'd688,  -14'd1149,  14'd1963,  
14'd1301,  -14'd50,  14'd361,  14'd749,  -14'd1124,  14'd603,  14'd384,  -14'd433,  -14'd595,  14'd1150,  14'd1605,  14'd650,  -14'd385,  14'd361,  -14'd819,  -14'd125,  
-14'd829,  14'd296,  -14'd499,  14'd573,  -14'd175,  -14'd590,  14'd332,  14'd118,  14'd738,  -14'd418,  14'd175,  14'd2153,  -14'd356,  -14'd769,  14'd235,  14'd241,  
14'd13,  -14'd787,  -14'd141,  14'd1178,  14'd806,  14'd2016,  -14'd640,  14'd1044,  14'd1088,  -14'd1103,  14'd1101,  -14'd1447,  14'd615,  14'd303,  14'd1257,  14'd1360,  
-14'd1035,  -14'd244,  14'd862,  14'd2336,  -14'd35,  -14'd509,  14'd987,  -14'd1421,  14'd1343,  -14'd2094,  -14'd1357,  -14'd232,  14'd358,  14'd614,  14'd657,  -14'd565,  
14'd944,  14'd893,  -14'd1674,  -14'd190,  -14'd698,  14'd303,  14'd83,  -14'd314,  14'd427,  14'd1937,  -14'd153,  -14'd1680,  14'd225,  14'd303,  -14'd1056,  -14'd134,  
14'd602,  14'd1310,  -14'd98,  -14'd587,  14'd155,  -14'd1528,  14'd147,  -14'd1291,  
14'd863,  14'd431,  14'd1542,  14'd419,  -14'd528,  14'd307,  14'd1028,  14'd2360,  -14'd173,  14'd1288,  -14'd1203,  -14'd441,  -14'd514,  -14'd119,  -14'd990,  -14'd1862,  
-14'd1512,  14'd868,  14'd467,  -14'd543,  -14'd695,  -14'd818,  -14'd714,  14'd913,  -14'd503,  -14'd379,  14'd1198,  14'd124,  -14'd957,  14'd819,  -14'd383,  -14'd232,  
-14'd569,  -14'd190,  -14'd569,  14'd1188,  14'd354,  14'd43,  14'd914,  14'd157,  14'd1300,  -14'd299,  14'd326,  -14'd178,  14'd480,  -14'd444,  -14'd317,  14'd955,  
14'd913,  14'd1552,  14'd63,  -14'd2244,  -14'd1579,  -14'd768,  14'd494,  -14'd87,  14'd778,  -14'd319,  14'd1604,  14'd219,  14'd447,  14'd573,  14'd986,  14'd838,  
-14'd1189,  14'd442,  -14'd1481,  -14'd1522,  -14'd912,  -14'd917,  -14'd1590,  14'd444,  -14'd1498,  14'd300,  14'd820,  14'd35,  14'd1804,  -14'd433,  14'd259,  14'd489,  
14'd947,  -14'd513,  14'd552,  14'd65,  14'd573,  14'd954,  14'd769,  14'd1218,  14'd704,  -14'd414,  14'd1306,  -14'd1412,  -14'd159,  14'd1349,  14'd505,  -14'd376,  
-14'd346,  -14'd182,  14'd862,  -14'd259,  14'd1288,  14'd250,  14'd1374,  14'd950,  14'd127,  -14'd711,  -14'd674,  -14'd1541,  -14'd332,  -14'd2095,  -14'd560,  -14'd587,  
14'd545,  -14'd170,  -14'd822,  14'd391,  14'd319,  -14'd1004,  14'd323,  14'd997,  
-14'd533,  14'd672,  14'd837,  -14'd190,  -14'd111,  -14'd469,  -14'd213,  14'd672,  -14'd118,  14'd1660,  14'd830,  -14'd1320,  14'd172,  -14'd908,  14'd453,  -14'd2675,  
-14'd265,  14'd1048,  14'd130,  -14'd743,  14'd100,  -14'd82,  14'd540,  14'd768,  -14'd654,  -14'd368,  -14'd990,  -14'd2655,  -14'd72,  -14'd789,  14'd978,  14'd749,  
-14'd562,  14'd954,  -14'd556,  14'd775,  14'd149,  -14'd2930,  -14'd882,  -14'd696,  -14'd181,  -14'd1284,  14'd980,  -14'd155,  14'd1047,  14'd1619,  -14'd56,  14'd645,  
14'd535,  14'd880,  14'd645,  -14'd609,  -14'd1392,  -14'd1384,  -14'd1461,  14'd306,  -14'd415,  14'd1242,  14'd847,  -14'd239,  -14'd1761,  -14'd528,  -14'd1074,  14'd94,  
14'd660,  14'd826,  -14'd67,  14'd662,  -14'd613,  14'd164,  14'd1377,  -14'd390,  -14'd1251,  -14'd1620,  14'd386,  14'd771,  14'd903,  14'd1388,  14'd80,  -14'd516,  
14'd215,  14'd265,  14'd1235,  14'd1161,  14'd423,  -14'd13,  -14'd1852,  -14'd1032,  14'd256,  -14'd1236,  14'd681,  -14'd255,  -14'd122,  14'd1274,  14'd62,  -14'd1314,  
14'd1690,  -14'd400,  14'd1385,  -14'd614,  14'd55,  14'd45,  -14'd340,  14'd1253,  14'd317,  14'd12,  -14'd857,  -14'd2660,  -14'd141,  -14'd632,  -14'd2259,  14'd1217,  
-14'd714,  14'd1231,  -14'd1927,  -14'd439,  -14'd1090,  -14'd604,  14'd860,  14'd791,  
-14'd73,  14'd1019,  14'd403,  14'd57,  14'd911,  -14'd312,  -14'd449,  14'd2341,  14'd1295,  -14'd528,  14'd37,  -14'd208,  14'd1,  14'd137,  14'd1636,  14'd393,  
14'd78,  -14'd524,  -14'd670,  14'd1389,  14'd1405,  14'd396,  14'd1064,  14'd166,  14'd646,  -14'd174,  -14'd169,  -14'd143,  14'd1106,  14'd1611,  14'd1027,  14'd1199,  
-14'd771,  -14'd294,  -14'd337,  14'd891,  -14'd1382,  14'd828,  14'd59,  14'd1455,  -14'd1184,  -14'd561,  14'd1622,  14'd461,  -14'd11,  14'd501,  14'd36,  14'd1275,  
-14'd1474,  14'd226,  -14'd18,  14'd1165,  -14'd791,  14'd53,  -14'd769,  -14'd65,  14'd461,  -14'd2216,  -14'd336,  14'd1140,  -14'd975,  14'd1759,  14'd619,  14'd207,  
-14'd869,  -14'd552,  -14'd109,  14'd592,  14'd138,  -14'd222,  -14'd360,  -14'd534,  14'd661,  -14'd170,  -14'd51,  14'd59,  14'd594,  -14'd5,  -14'd371,  -14'd1077,  
-14'd1098,  14'd341,  14'd953,  14'd114,  -14'd156,  14'd266,  -14'd269,  -14'd523,  14'd780,  -14'd544,  14'd512,  14'd539,  -14'd26,  14'd13,  14'd450,  -14'd303,  
14'd377,  14'd1047,  -14'd2620,  14'd477,  -14'd27,  -14'd687,  -14'd1431,  -14'd948,  14'd63,  14'd555,  14'd76,  -14'd251,  -14'd479,  -14'd1192,  -14'd1512,  -14'd18,  
14'd1003,  14'd2152,  -14'd379,  14'd329,  -14'd862,  14'd224,  14'd549,  -14'd1175,  
-14'd810,  14'd587,  -14'd1377,  14'd274,  -14'd115,  14'd257,  -14'd953,  -14'd2685,  -14'd2035,  -14'd1273,  -14'd294,  -14'd1202,  -14'd1748,  -14'd168,  -14'd794,  -14'd101,  
-14'd1027,  -14'd890,  -14'd77,  -14'd743,  -14'd985,  -14'd379,  -14'd116,  14'd397,  -14'd131,  -14'd817,  -14'd1033,  -14'd105,  -14'd422,  -14'd872,  -14'd550,  -14'd25,  
-14'd239,  14'd1184,  14'd975,  -14'd718,  14'd610,  -14'd361,  -14'd796,  14'd929,  -14'd701,  14'd107,  14'd259,  14'd949,  14'd521,  -14'd178,  -14'd556,  -14'd1170,  
-14'd389,  -14'd254,  14'd558,  14'd625,  14'd288,  -14'd976,  14'd626,  -14'd710,  -14'd503,  -14'd1548,  -14'd732,  -14'd1339,  -14'd1698,  -14'd538,  14'd73,  -14'd89,  
-14'd588,  14'd341,  14'd572,  14'd1146,  14'd5,  -14'd389,  14'd1846,  -14'd1336,  14'd303,  -14'd831,  14'd997,  -14'd576,  -14'd805,  -14'd1568,  -14'd1476,  -14'd939,  
14'd12,  -14'd766,  14'd9,  -14'd988,  -14'd999,  -14'd1042,  14'd661,  14'd294,  -14'd1003,  -14'd440,  14'd484,  14'd447,  14'd366,  -14'd156,  14'd516,  -14'd785,  
-14'd1652,  -14'd452,  14'd1106,  14'd1193,  14'd972,  -14'd86,  -14'd1324,  -14'd1840,  14'd152,  -14'd1233,  -14'd575,  -14'd1120,  14'd559,  -14'd522,  -14'd155,  -14'd1098,  
-14'd43,  14'd261,  -14'd28,  14'd76,  -14'd370,  14'd123,  -14'd0,  -14'd1203,  
-14'd61,  14'd962,  14'd357,  -14'd952,  14'd66,  -14'd719,  14'd438,  -14'd350,  14'd249,  14'd55,  14'd995,  -14'd706,  -14'd862,  -14'd719,  -14'd237,  -14'd20,  
14'd1824,  14'd687,  -14'd64,  14'd1334,  -14'd578,  14'd793,  -14'd235,  -14'd2893,  14'd242,  -14'd666,  14'd705,  14'd1078,  -14'd245,  -14'd190,  14'd1179,  -14'd883,  
14'd284,  14'd534,  -14'd1051,  14'd1060,  -14'd995,  14'd987,  -14'd186,  14'd157,  -14'd1628,  14'd1168,  -14'd148,  14'd830,  -14'd1179,  14'd1352,  14'd66,  14'd145,  
14'd568,  14'd1347,  14'd1397,  -14'd329,  -14'd182,  14'd229,  14'd1751,  -14'd899,  14'd982,  -14'd1244,  -14'd756,  -14'd1942,  14'd219,  14'd395,  14'd471,  -14'd1304,  
-14'd962,  14'd1392,  14'd271,  14'd427,  -14'd220,  -14'd1510,  14'd388,  14'd469,  14'd1700,  -14'd696,  14'd299,  -14'd940,  -14'd2160,  -14'd300,  -14'd1688,  -14'd412,  
14'd596,  -14'd40,  14'd546,  -14'd218,  14'd1865,  14'd1372,  14'd586,  -14'd593,  -14'd1063,  -14'd1664,  14'd15,  14'd1000,  -14'd721,  14'd281,  14'd94,  -14'd692,  
14'd415,  -14'd277,  -14'd585,  14'd38,  14'd1467,  14'd578,  -14'd891,  -14'd815,  14'd1492,  -14'd660,  14'd140,  14'd598,  -14'd599,  14'd2550,  -14'd796,  -14'd744,  
14'd245,  14'd1298,  -14'd31,  -14'd1365,  -14'd744,  14'd885,  14'd262,  -14'd63,  
-14'd1431,  14'd89,  -14'd1234,  14'd653,  14'd453,  14'd1160,  14'd183,  14'd976,  -14'd1660,  14'd1485,  -14'd2036,  14'd766,  14'd296,  14'd1459,  14'd732,  -14'd1715,  
14'd1486,  14'd1331,  -14'd505,  -14'd834,  -14'd757,  14'd247,  14'd635,  14'd798,  -14'd274,  -14'd13,  -14'd368,  14'd586,  14'd2229,  14'd952,  14'd2672,  14'd279,  
-14'd438,  14'd1423,  14'd367,  14'd393,  14'd229,  -14'd1150,  -14'd193,  -14'd161,  14'd556,  -14'd893,  -14'd1312,  -14'd1266,  -14'd212,  14'd288,  -14'd533,  14'd687,  
-14'd1286,  -14'd349,  -14'd41,  -14'd327,  14'd385,  -14'd1130,  -14'd2228,  14'd642,  14'd262,  14'd1362,  14'd451,  14'd547,  -14'd450,  14'd686,  -14'd147,  -14'd232,  
-14'd361,  14'd645,  -14'd905,  -14'd726,  -14'd57,  -14'd1135,  -14'd239,  14'd686,  -14'd835,  -14'd290,  -14'd169,  14'd758,  -14'd449,  14'd862,  -14'd1053,  14'd644,  
14'd762,  14'd604,  14'd710,  14'd812,  -14'd327,  -14'd952,  -14'd201,  14'd820,  14'd655,  -14'd796,  -14'd1824,  14'd1405,  -14'd1175,  -14'd1,  14'd1534,  14'd297,  
14'd782,  -14'd699,  14'd70,  -14'd755,  14'd748,  14'd49,  -14'd1011,  -14'd1714,  -14'd146,  14'd368,  14'd233,  14'd568,  -14'd459,  -14'd845,  14'd314,  -14'd1102,  
14'd2133,  -14'd538,  -14'd1178,  14'd40,  14'd872,  -14'd1024,  14'd232,  -14'd900,  
14'd1237,  -14'd47,  14'd1409,  14'd207,  -14'd746,  14'd1328,  -14'd1400,  14'd845,  -14'd1094,  -14'd1304,  14'd197,  14'd308,  -14'd879,  14'd172,  14'd431,  -14'd247,  
14'd844,  -14'd720,  14'd782,  14'd791,  -14'd752,  -14'd622,  14'd189,  -14'd62,  -14'd246,  -14'd88,  14'd1492,  14'd1228,  -14'd1559,  -14'd357,  -14'd22,  14'd12,  
-14'd258,  -14'd612,  14'd73,  14'd932,  14'd1134,  -14'd814,  14'd255,  -14'd1233,  14'd1255,  14'd1622,  14'd1859,  -14'd546,  -14'd303,  -14'd1271,  14'd278,  -14'd1028,  
14'd62,  14'd233,  14'd489,  14'd1055,  14'd230,  -14'd96,  14'd597,  -14'd1424,  -14'd1418,  14'd71,  -14'd775,  -14'd1572,  14'd206,  -14'd517,  14'd1107,  14'd97,  
14'd167,  14'd1356,  14'd509,  -14'd69,  14'd767,  14'd1579,  14'd577,  14'd131,  14'd1058,  -14'd538,  -14'd473,  14'd348,  -14'd244,  -14'd1386,  -14'd1974,  -14'd1259,  
-14'd668,  14'd689,  -14'd285,  -14'd1106,  14'd1162,  14'd531,  14'd709,  14'd60,  14'd1126,  14'd1757,  14'd568,  14'd398,  -14'd602,  14'd1517,  -14'd274,  14'd1793,  
-14'd485,  -14'd1469,  14'd593,  -14'd248,  14'd414,  -14'd933,  14'd356,  14'd2066,  14'd379,  -14'd26,  -14'd404,  14'd1713,  14'd1115,  14'd942,  14'd2077,  14'd396,  
-14'd384,  -14'd141,  14'd1732,  14'd55,  14'd86,  -14'd1304,  -14'd1688,  14'd717,  
-14'd1589,  14'd740,  -14'd74,  -14'd712,  -14'd671,  14'd1310,  14'd625,  -14'd445,  14'd323,  -14'd340,  -14'd1138,  -14'd509,  -14'd1007,  14'd317,  -14'd468,  14'd37,  
-14'd144,  14'd1266,  14'd721,  14'd232,  14'd1159,  -14'd1210,  -14'd602,  14'd901,  -14'd861,  14'd336,  -14'd405,  -14'd1259,  -14'd1164,  -14'd150,  14'd77,  14'd965,  
-14'd680,  14'd459,  14'd142,  14'd1,  -14'd204,  -14'd1177,  -14'd109,  -14'd851,  14'd372,  14'd81,  -14'd215,  -14'd232,  -14'd377,  -14'd223,  14'd497,  -14'd603,  
14'd223,  -14'd877,  14'd1482,  -14'd320,  -14'd471,  -14'd1554,  14'd488,  14'd628,  -14'd249,  -14'd798,  14'd844,  -14'd1752,  -14'd186,  -14'd206,  -14'd737,  14'd166,  
14'd267,  -14'd368,  -14'd151,  -14'd520,  14'd447,  14'd183,  14'd366,  14'd812,  -14'd129,  14'd1061,  -14'd32,  -14'd1169,  -14'd284,  -14'd89,  -14'd1109,  14'd707,  
14'd296,  -14'd536,  -14'd860,  -14'd442,  -14'd370,  -14'd385,  -14'd330,  14'd319,  14'd5,  -14'd348,  -14'd673,  -14'd958,  -14'd659,  -14'd823,  -14'd50,  14'd109,  
14'd416,  -14'd984,  -14'd1407,  14'd1006,  -14'd687,  -14'd674,  -14'd690,  -14'd1609,  -14'd178,  14'd110,  -14'd182,  -14'd554,  -14'd153,  -14'd347,  -14'd689,  14'd1331,  
14'd557,  14'd898,  14'd894,  14'd430,  -14'd721,  14'd244,  14'd432,  -14'd790,  
14'd1667,  14'd551,  -14'd1556,  -14'd696,  14'd134,  -14'd893,  -14'd57,  14'd717,  -14'd444,  -14'd1101,  -14'd2251,  -14'd910,  14'd1035,  -14'd789,  14'd708,  -14'd8,  
14'd1643,  -14'd284,  14'd322,  14'd2113,  -14'd1257,  14'd716,  14'd1554,  14'd2315,  14'd63,  -14'd572,  14'd316,  -14'd665,  14'd194,  14'd112,  14'd1628,  -14'd151,  
14'd69,  -14'd866,  -14'd1020,  14'd994,  -14'd877,  14'd1434,  14'd1887,  -14'd660,  14'd874,  14'd20,  14'd566,  14'd234,  -14'd951,  -14'd1287,  -14'd412,  14'd250,  
14'd347,  -14'd65,  -14'd818,  14'd1075,  14'd718,  -14'd1265,  -14'd208,  14'd111,  14'd170,  14'd944,  -14'd883,  -14'd1529,  -14'd894,  -14'd336,  -14'd1739,  14'd249,  
14'd1428,  -14'd521,  14'd623,  14'd2372,  -14'd1450,  14'd356,  -14'd247,  14'd615,  14'd385,  -14'd232,  -14'd660,  -14'd774,  14'd86,  -14'd170,  14'd564,  14'd94,  
-14'd184,  14'd1189,  -14'd216,  14'd822,  14'd686,  -14'd554,  14'd1195,  -14'd323,  14'd1497,  14'd1130,  -14'd335,  14'd192,  14'd424,  14'd1301,  -14'd982,  14'd823,  
14'd824,  -14'd767,  -14'd5,  14'd1648,  14'd244,  -14'd56,  14'd674,  14'd1863,  -14'd237,  14'd23,  14'd1008,  14'd566,  14'd1454,  14'd1013,  14'd1689,  14'd137,  
-14'd135,  14'd1056,  14'd509,  14'd1010,  14'd1377,  14'd1307,  14'd671,  14'd96,  
14'd541,  14'd718,  -14'd1658,  14'd674,  14'd454,  14'd778,  14'd66,  14'd809,  14'd552,  14'd275,  -14'd1518,  -14'd958,  14'd1250,  -14'd1488,  14'd93,  14'd885,  
14'd1055,  -14'd723,  14'd147,  -14'd1153,  14'd294,  14'd111,  14'd1283,  14'd944,  14'd1351,  -14'd892,  -14'd544,  14'd324,  14'd941,  -14'd392,  14'd837,  14'd526,  
14'd504,  14'd892,  14'd1046,  -14'd132,  -14'd1525,  -14'd738,  -14'd222,  14'd430,  -14'd230,  -14'd535,  14'd375,  -14'd968,  14'd1882,  14'd885,  -14'd601,  -14'd369,  
14'd504,  -14'd148,  14'd615,  -14'd284,  -14'd1168,  -14'd1097,  -14'd583,  -14'd779,  14'd1979,  -14'd519,  -14'd1156,  14'd385,  -14'd9,  14'd1067,  -14'd436,  14'd23,  
-14'd1273,  14'd2205,  14'd680,  -14'd225,  14'd107,  -14'd1164,  14'd612,  -14'd1321,  14'd543,  14'd63,  14'd1340,  14'd355,  14'd1516,  -14'd25,  14'd1185,  -14'd352,  
14'd45,  14'd1702,  14'd292,  14'd306,  -14'd1494,  -14'd578,  14'd635,  -14'd551,  -14'd858,  -14'd688,  -14'd49,  -14'd308,  -14'd292,  -14'd194,  -14'd378,  14'd973,  
-14'd117,  14'd518,  -14'd11,  -14'd665,  14'd967,  14'd514,  14'd671,  -14'd1445,  -14'd1302,  14'd1063,  14'd1790,  -14'd2097,  14'd805,  14'd587,  -14'd112,  14'd887,  
-14'd428,  -14'd681,  -14'd54,  14'd904,  -14'd398,  -14'd1597,  -14'd178,  14'd102,  
14'd402,  -14'd473,  14'd79,  14'd469,  -14'd1139,  -14'd569,  -14'd245,  -14'd510,  14'd60,  -14'd228,  -14'd1781,  14'd1740,  14'd1560,  14'd693,  14'd878,  14'd760,  
-14'd68,  14'd1071,  -14'd30,  -14'd411,  14'd293,  -14'd632,  14'd1058,  14'd849,  -14'd720,  14'd383,  -14'd248,  -14'd749,  14'd751,  14'd681,  -14'd1300,  14'd1771,  
14'd176,  14'd373,  14'd401,  14'd930,  14'd1626,  -14'd1324,  -14'd506,  14'd278,  14'd1573,  14'd859,  -14'd1077,  14'd473,  -14'd1852,  -14'd285,  14'd164,  -14'd1896,  
14'd425,  -14'd1868,  14'd825,  14'd1991,  -14'd1570,  14'd1258,  14'd1105,  -14'd583,  14'd119,  14'd170,  -14'd761,  -14'd768,  14'd621,  -14'd544,  -14'd1206,  -14'd816,  
-14'd369,  -14'd87,  14'd813,  -14'd174,  -14'd269,  -14'd1098,  -14'd532,  14'd1135,  14'd444,  14'd503,  14'd1070,  14'd304,  14'd1037,  -14'd303,  14'd1151,  14'd317,  
-14'd546,  -14'd1494,  -14'd71,  -14'd1690,  -14'd438,  14'd790,  14'd1185,  14'd854,  14'd1198,  -14'd17,  14'd776,  14'd805,  -14'd1347,  14'd1490,  14'd160,  -14'd243,  
14'd254,  -14'd319,  14'd994,  -14'd1211,  -14'd291,  -14'd86,  -14'd36,  -14'd1145,  14'd938,  14'd169,  14'd2455,  14'd128,  -14'd190,  14'd1750,  -14'd714,  14'd1961,  
14'd1598,  -14'd1052,  14'd855,  14'd1085,  14'd465,  -14'd758,  -14'd449,  -14'd283,  
14'd249,  14'd316,  14'd1331,  14'd226,  14'd610,  14'd208,  14'd1275,  14'd239,  14'd287,  -14'd174,  14'd662,  -14'd93,  14'd317,  14'd138,  -14'd954,  -14'd41,  
14'd333,  14'd541,  14'd1232,  14'd660,  14'd973,  14'd306,  -14'd1014,  -14'd1432,  14'd348,  14'd20,  -14'd850,  14'd163,  14'd440,  14'd11,  -14'd1123,  -14'd641,  
14'd378,  14'd1435,  -14'd456,  -14'd803,  14'd1003,  -14'd182,  -14'd1149,  -14'd860,  -14'd495,  -14'd539,  14'd2403,  14'd1771,  -14'd208,  14'd461,  14'd410,  -14'd909,  
-14'd109,  14'd1719,  14'd500,  14'd1306,  -14'd1143,  14'd875,  -14'd1103,  -14'd209,  14'd121,  -14'd5,  -14'd1167,  -14'd712,  14'd983,  -14'd439,  14'd2061,  -14'd1653,  
-14'd1546,  14'd671,  14'd724,  -14'd554,  14'd378,  14'd469,  -14'd287,  -14'd65,  14'd1583,  -14'd772,  -14'd9,  14'd1717,  -14'd74,  14'd843,  -14'd115,  -14'd1054,  
14'd22,  -14'd289,  14'd2108,  14'd1454,  14'd292,  14'd194,  14'd414,  -14'd1282,  -14'd12,  14'd393,  14'd334,  -14'd558,  -14'd727,  14'd1197,  -14'd454,  -14'd614,  
14'd478,  -14'd951,  14'd1488,  14'd1038,  14'd1421,  14'd1362,  -14'd259,  -14'd248,  -14'd880,  14'd1059,  -14'd713,  -14'd684,  -14'd57,  -14'd436,  -14'd1324,  14'd1847,  
14'd415,  -14'd94,  14'd920,  -14'd345,  -14'd384,  -14'd368,  -14'd583,  -14'd176,  
14'd859,  -14'd33,  -14'd1642,  14'd561,  -14'd1173,  -14'd429,  14'd927,  -14'd18,  14'd951,  14'd1522,  14'd627,  14'd528,  -14'd324,  14'd1892,  14'd274,  -14'd2541,  
-14'd2052,  -14'd67,  -14'd1552,  14'd1518,  14'd271,  14'd96,  14'd645,  -14'd1007,  14'd687,  -14'd323,  14'd1867,  -14'd206,  14'd195,  14'd2309,  14'd496,  14'd767,  
-14'd705,  -14'd1294,  -14'd1510,  -14'd1401,  14'd1029,  -14'd434,  -14'd57,  -14'd301,  14'd945,  14'd411,  -14'd1653,  -14'd1215,  14'd388,  14'd1255,  -14'd1042,  14'd1614,  
14'd135,  -14'd1877,  -14'd190,  -14'd616,  -14'd31,  -14'd1349,  -14'd159,  -14'd138,  14'd453,  14'd2194,  14'd88,  -14'd525,  14'd1065,  14'd257,  -14'd896,  -14'd1377,  
14'd1267,  -14'd500,  14'd861,  14'd966,  -14'd467,  -14'd438,  -14'd1950,  14'd212,  -14'd219,  14'd668,  -14'd518,  14'd1549,  14'd1290,  -14'd268,  14'd410,  -14'd834,  
-14'd556,  -14'd647,  -14'd270,  14'd918,  14'd194,  14'd121,  -14'd1890,  14'd714,  -14'd470,  14'd880,  -14'd914,  14'd1132,  14'd702,  -14'd354,  -14'd1005,  -14'd1055,  
-14'd497,  -14'd574,  -14'd146,  -14'd1502,  14'd915,  -14'd2474,  14'd1305,  14'd2453,  14'd549,  -14'd158,  -14'd1059,  14'd430,  14'd164,  14'd1073,  14'd1428,  -14'd1167,  
-14'd763,  14'd1158,  14'd1521,  14'd609,  14'd121,  -14'd1466,  -14'd961,  -14'd782,  
14'd50,  14'd218,  -14'd767,  14'd224,  14'd744,  -14'd181,  -14'd1955,  -14'd838,  14'd599,  -14'd31,  14'd649,  -14'd395,  -14'd501,  -14'd303,  -14'd390,  -14'd1219,  
-14'd1514,  14'd743,  -14'd443,  14'd79,  -14'd796,  -14'd553,  14'd130,  14'd474,  14'd468,  -14'd794,  14'd87,  -14'd442,  14'd64,  -14'd423,  -14'd71,  -14'd1077,  
14'd653,  -14'd1451,  14'd915,  14'd27,  -14'd88,  -14'd1167,  14'd173,  -14'd1884,  14'd205,  -14'd120,  14'd1274,  -14'd1349,  -14'd1769,  14'd699,  -14'd451,  -14'd311,  
-14'd757,  14'd523,  14'd63,  -14'd905,  -14'd46,  -14'd1042,  -14'd713,  -14'd382,  -14'd686,  14'd211,  -14'd1483,  -14'd1315,  -14'd647,  -14'd1437,  -14'd219,  -14'd1123,  
-14'd84,  -14'd688,  14'd132,  -14'd1488,  14'd66,  -14'd590,  -14'd1894,  -14'd808,  -14'd206,  -14'd1428,  -14'd499,  -14'd485,  14'd751,  14'd654,  -14'd9,  14'd728,  
-14'd1375,  -14'd656,  -14'd1906,  -14'd14,  -14'd1331,  -14'd928,  -14'd1990,  -14'd358,  -14'd170,  14'd116,  -14'd12,  -14'd227,  -14'd994,  -14'd1306,  -14'd274,  14'd831,  
-14'd1097,  -14'd886,  -14'd617,  14'd41,  -14'd1665,  14'd148,  14'd1113,  -14'd618,  14'd201,  -14'd1083,  -14'd27,  -14'd533,  -14'd1107,  -14'd1080,  -14'd446,  -14'd301,  
-14'd480,  14'd332,  -14'd90,  -14'd208,  14'd354,  14'd279,  -14'd612,  14'd896,  
14'd2370,  -14'd258,  14'd1422,  -14'd401,  14'd2031,  -14'd359,  -14'd477,  14'd659,  -14'd1981,  -14'd228,  -14'd333,  14'd514,  -14'd1633,  14'd1849,  -14'd157,  -14'd1232,  
14'd1955,  14'd382,  -14'd168,  14'd339,  14'd260,  -14'd515,  -14'd998,  14'd776,  14'd37,  14'd1791,  14'd353,  -14'd1562,  -14'd1031,  14'd1114,  -14'd224,  14'd832,  
-14'd243,  14'd221,  14'd160,  -14'd581,  -14'd40,  14'd1231,  14'd280,  14'd253,  14'd1069,  14'd673,  14'd1769,  -14'd468,  14'd161,  14'd203,  14'd54,  -14'd1797,  
14'd559,  -14'd233,  14'd1573,  14'd1730,  -14'd3,  14'd1604,  14'd477,  -14'd115,  14'd71,  -14'd314,  -14'd302,  -14'd147,  14'd982,  14'd237,  -14'd1153,  -14'd1937,  
14'd265,  -14'd381,  -14'd294,  -14'd1672,  -14'd524,  14'd237,  14'd656,  14'd778,  14'd1142,  14'd411,  14'd1131,  -14'd853,  14'd482,  14'd924,  14'd1352,  14'd660,  
-14'd889,  14'd880,  14'd39,  -14'd24,  -14'd111,  -14'd866,  -14'd1418,  -14'd762,  -14'd1429,  -14'd103,  14'd1780,  -14'd56,  -14'd405,  14'd301,  14'd752,  -14'd1883,  
-14'd1008,  -14'd1166,  14'd227,  14'd745,  14'd1374,  14'd1197,  14'd392,  -14'd233,  14'd740,  14'd383,  14'd618,  14'd42,  14'd1208,  -14'd2037,  14'd54,  14'd797,  
-14'd605,  14'd1864,  -14'd857,  14'd1051,  14'd40,  -14'd444,  -14'd458,  14'd260,  
-14'd1028,  -14'd640,  -14'd9,  -14'd921,  14'd386,  -14'd528,  14'd843,  14'd68,  14'd651,  -14'd604,  -14'd939,  14'd187,  -14'd126,  -14'd160,  -14'd596,  14'd2,  
-14'd847,  14'd605,  14'd918,  -14'd1041,  -14'd679,  14'd515,  -14'd379,  14'd1107,  -14'd395,  14'd886,  14'd1285,  14'd514,  -14'd173,  14'd1054,  -14'd858,  -14'd951,  
14'd231,  -14'd391,  14'd392,  -14'd291,  -14'd663,  14'd896,  14'd1288,  -14'd284,  -14'd454,  14'd451,  -14'd949,  14'd1421,  -14'd104,  -14'd795,  -14'd142,  14'd1329,  
14'd459,  14'd145,  -14'd600,  -14'd2175,  14'd165,  -14'd244,  -14'd259,  14'd155,  14'd1224,  -14'd1243,  -14'd1481,  -14'd1255,  14'd735,  -14'd209,  -14'd2280,  14'd202,  
14'd648,  -14'd1419,  14'd7,  14'd1392,  14'd1573,  14'd105,  14'd106,  14'd1010,  14'd759,  14'd254,  14'd181,  14'd947,  -14'd1870,  -14'd112,  14'd804,  -14'd793,  
14'd1221,  14'd44,  -14'd19,  14'd1019,  14'd183,  -14'd1513,  14'd777,  14'd1411,  -14'd540,  14'd714,  14'd1803,  14'd663,  -14'd89,  14'd27,  -14'd614,  14'd859,  
-14'd719,  -14'd169,  -14'd360,  14'd363,  -14'd602,  14'd774,  -14'd718,  14'd2521,  14'd138,  14'd862,  -14'd277,  -14'd740,  14'd409,  -14'd1351,  -14'd122,  14'd697,  
-14'd999,  14'd332,  -14'd1207,  -14'd875,  14'd235,  14'd1099,  14'd39,  14'd737,  
-14'd57,  14'd63,  -14'd1110,  -14'd1500,  14'd1093,  14'd1975,  14'd103,  -14'd937,  -14'd517,  -14'd1257,  14'd272,  14'd609,  14'd626,  14'd1391,  14'd545,  14'd1145,  
14'd809,  14'd123,  -14'd1532,  -14'd1535,  14'd258,  -14'd277,  -14'd807,  14'd757,  14'd1140,  -14'd1735,  -14'd48,  -14'd1056,  -14'd793,  14'd951,  14'd518,  14'd84,  
-14'd463,  14'd486,  -14'd819,  14'd135,  14'd71,  14'd377,  -14'd1141,  14'd373,  -14'd939,  14'd1249,  -14'd395,  -14'd138,  -14'd295,  14'd346,  -14'd587,  -14'd1285,  
14'd869,  14'd521,  14'd396,  -14'd2301,  -14'd9,  -14'd715,  14'd911,  -14'd514,  -14'd93,  -14'd122,  -14'd928,  -14'd966,  -14'd1355,  14'd661,  -14'd497,  14'd594,  
14'd1176,  -14'd39,  -14'd718,  14'd168,  14'd505,  -14'd2571,  14'd1037,  14'd472,  14'd1351,  -14'd1981,  14'd857,  -14'd243,  14'd222,  -14'd340,  14'd230,  -14'd1184,  
14'd81,  14'd517,  14'd899,  -14'd1362,  14'd632,  14'd898,  14'd347,  -14'd316,  14'd1527,  14'd300,  14'd648,  14'd677,  14'd636,  -14'd527,  -14'd692,  14'd294,  
-14'd345,  -14'd35,  14'd1420,  14'd1319,  14'd788,  14'd204,  -14'd334,  -14'd689,  -14'd153,  14'd975,  14'd1442,  -14'd422,  -14'd999,  -14'd427,  14'd127,  -14'd180,  
14'd65,  14'd160,  -14'd488,  -14'd173,  -14'd534,  -14'd882,  14'd272,  14'd1134,  
14'd22,  -14'd30,  14'd86,  -14'd277,  14'd729,  -14'd464,  -14'd1890,  14'd1132,  -14'd2466,  -14'd308,  -14'd1520,  -14'd781,  14'd534,  14'd927,  14'd717,  14'd85,  
-14'd972,  14'd1463,  -14'd1750,  -14'd348,  -14'd1094,  -14'd972,  14'd360,  14'd1985,  -14'd31,  14'd1010,  -14'd141,  -14'd1754,  14'd913,  14'd1372,  -14'd1373,  14'd1932,  
-14'd1542,  -14'd16,  14'd511,  14'd600,  14'd2243,  14'd1074,  14'd234,  -14'd562,  14'd457,  14'd247,  -14'd344,  -14'd1156,  14'd70,  -14'd1384,  -14'd894,  -14'd2506,  
14'd863,  -14'd725,  -14'd1510,  14'd460,  14'd782,  14'd168,  -14'd1620,  14'd20,  -14'd733,  -14'd387,  14'd834,  14'd195,  -14'd333,  14'd1070,  -14'd784,  14'd53,  
14'd1185,  -14'd384,  -14'd528,  14'd266,  -14'd155,  -14'd1186,  14'd601,  -14'd223,  14'd412,  -14'd988,  14'd734,  -14'd223,  -14'd2108,  14'd564,  14'd187,  -14'd878,  
-14'd781,  14'd632,  -14'd1932,  -14'd78,  -14'd706,  14'd50,  -14'd612,  -14'd551,  -14'd54,  -14'd186,  -14'd206,  -14'd684,  -14'd151,  -14'd920,  -14'd771,  14'd770,  
14'd423,  -14'd628,  -14'd424,  -14'd2449,  14'd93,  -14'd27,  -14'd109,  14'd31,  -14'd670,  14'd1039,  14'd196,  -14'd1830,  -14'd671,  14'd1730,  14'd422,  14'd1618,  
-14'd767,  -14'd1063,  14'd850,  14'd213,  14'd432,  14'd320,  14'd1793,  14'd389,  
-14'd788,  -14'd1266,  -14'd620,  -14'd402,  14'd556,  14'd42,  14'd152,  14'd68,  -14'd149,  14'd1380,  -14'd524,  14'd1169,  14'd148,  14'd345,  -14'd1004,  14'd332,  
-14'd81,  -14'd128,  14'd13,  -14'd100,  -14'd627,  -14'd871,  -14'd949,  14'd806,  -14'd501,  14'd139,  14'd308,  14'd1106,  -14'd162,  -14'd691,  -14'd1367,  14'd871,  
-14'd1826,  -14'd2,  14'd1095,  -14'd192,  -14'd1418,  -14'd257,  14'd702,  14'd853,  14'd900,  -14'd992,  14'd1419,  14'd1404,  -14'd477,  -14'd229,  -14'd842,  14'd542,  
14'd44,  14'd54,  14'd459,  14'd28,  14'd458,  -14'd724,  -14'd223,  -14'd553,  -14'd901,  14'd795,  14'd1320,  14'd97,  14'd1097,  -14'd493,  14'd138,  -14'd1397,  
-14'd235,  14'd160,  14'd348,  14'd61,  14'd423,  -14'd441,  -14'd445,  14'd19,  -14'd609,  14'd2495,  14'd10,  14'd111,  14'd102,  -14'd37,  -14'd1403,  14'd1037,  
14'd15,  -14'd568,  -14'd1142,  -14'd902,  -14'd546,  -14'd152,  -14'd1531,  14'd1356,  -14'd147,  14'd801,  14'd1683,  14'd1165,  14'd637,  14'd795,  -14'd1020,  14'd1433,  
-14'd1167,  -14'd530,  14'd1997,  14'd448,  14'd395,  14'd747,  14'd646,  14'd587,  -14'd1600,  -14'd80,  -14'd38,  14'd1832,  14'd80,  14'd371,  14'd373,  14'd341,  
14'd489,  -14'd1057,  -14'd840,  14'd102,  14'd1535,  14'd1786,  -14'd354,  -14'd29,  
-14'd1175,  -14'd606,  -14'd441,  -14'd232,  14'd1374,  -14'd660,  14'd1161,  14'd978,  14'd2249,  -14'd578,  14'd885,  -14'd435,  14'd255,  14'd757,  14'd1707,  14'd417,  
14'd99,  -14'd940,  -14'd46,  -14'd611,  -14'd102,  -14'd273,  14'd573,  14'd843,  -14'd228,  14'd2169,  14'd154,  14'd1053,  14'd1,  14'd188,  -14'd624,  -14'd1424,  
14'd1827,  -14'd250,  14'd552,  14'd327,  -14'd1360,  14'd166,  -14'd457,  14'd191,  -14'd1020,  -14'd387,  14'd981,  14'd38,  14'd2086,  14'd480,  -14'd1198,  14'd878,  
14'd65,  14'd438,  14'd98,  14'd572,  -14'd1347,  14'd1155,  -14'd2196,  -14'd227,  14'd392,  -14'd1873,  14'd487,  -14'd149,  -14'd549,  14'd904,  14'd1608,  14'd1748,  
14'd565,  14'd750,  14'd504,  -14'd612,  14'd1131,  14'd319,  14'd902,  14'd91,  14'd873,  14'd617,  14'd83,  14'd315,  14'd719,  -14'd169,  -14'd849,  14'd154,  
-14'd1363,  -14'd59,  14'd1336,  14'd1947,  14'd661,  14'd1253,  14'd1,  -14'd1087,  -14'd687,  14'd355,  14'd1074,  -14'd516,  14'd1484,  14'd646,  -14'd502,  -14'd1039,  
-14'd598,  -14'd863,  -14'd627,  14'd2247,  -14'd979,  14'd1145,  14'd624,  -14'd444,  14'd978,  -14'd896,  -14'd355,  14'd976,  -14'd41,  -14'd1167,  -14'd714,  -14'd194,  
14'd785,  14'd1788,  -14'd1926,  14'd250,  -14'd598,  -14'd1010,  14'd463,  -14'd1020,  
-14'd44,  -14'd240,  -14'd1590,  14'd718,  -14'd503,  14'd630,  14'd652,  -14'd5,  -14'd101,  14'd241,  -14'd418,  14'd84,  -14'd209,  14'd83,  14'd809,  -14'd651,  
-14'd1416,  -14'd495,  14'd1539,  14'd265,  14'd121,  -14'd753,  -14'd324,  -14'd1202,  -14'd1166,  -14'd44,  14'd1278,  14'd783,  -14'd841,  14'd512,  -14'd564,  -14'd747,  
-14'd1993,  14'd1526,  -14'd665,  14'd153,  -14'd13,  14'd143,  -14'd478,  14'd145,  14'd1230,  -14'd1036,  -14'd1034,  14'd329,  14'd76,  14'd492,  14'd1651,  14'd1795,  
14'd1207,  -14'd1001,  14'd1811,  -14'd151,  14'd352,  14'd1246,  -14'd394,  14'd6,  -14'd209,  14'd1336,  14'd1180,  14'd329,  14'd785,  -14'd17,  14'd2618,  14'd109,  
-14'd904,  -14'd209,  14'd397,  -14'd116,  14'd382,  -14'd328,  14'd708,  -14'd141,  14'd138,  14'd185,  -14'd1466,  14'd1386,  14'd359,  -14'd1601,  -14'd738,  -14'd828,  
14'd331,  -14'd447,  14'd905,  -14'd920,  -14'd1437,  14'd1131,  -14'd605,  -14'd533,  14'd777,  14'd1755,  14'd385,  14'd1364,  -14'd1032,  14'd111,  14'd505,  14'd1417,  
-14'd94,  -14'd1012,  14'd2225,  -14'd766,  14'd430,  -14'd312,  -14'd142,  14'd1622,  -14'd1259,  -14'd384,  -14'd484,  14'd619,  14'd583,  14'd479,  14'd872,  -14'd414,  
14'd294,  -14'd479,  14'd1705,  -14'd89,  -14'd74,  14'd333,  14'd126,  -14'd152,  
14'd608,  -14'd1127,  14'd805,  -14'd458,  14'd445,  14'd141,  -14'd423,  -14'd116,  14'd505,  14'd118,  -14'd1196,  -14'd3,  14'd1327,  14'd39,  14'd1529,  -14'd77,  
14'd373,  14'd529,  -14'd671,  14'd1038,  14'd490,  -14'd165,  14'd1342,  14'd2118,  14'd275,  14'd1062,  -14'd1250,  14'd3,  14'd217,  -14'd602,  14'd794,  14'd402,  
-14'd353,  14'd583,  14'd712,  -14'd1068,  14'd679,  -14'd918,  14'd194,  14'd776,  -14'd470,  14'd399,  14'd389,  -14'd209,  14'd1575,  -14'd1132,  -14'd241,  -14'd1713,  
14'd647,  14'd1122,  -14'd579,  -14'd819,  14'd724,  -14'd635,  -14'd1577,  14'd941,  14'd262,  14'd464,  -14'd372,  14'd1037,  14'd291,  14'd512,  -14'd1984,  14'd626,  
14'd1450,  -14'd76,  14'd649,  14'd402,  14'd1758,  14'd701,  -14'd875,  -14'd295,  -14'd688,  -14'd857,  14'd1064,  -14'd189,  14'd1321,  -14'd682,  14'd782,  -14'd186,  
14'd466,  14'd1848,  -14'd1572,  14'd1064,  -14'd2242,  -14'd1204,  14'd1238,  14'd1947,  -14'd117,  14'd94,  -14'd1111,  14'd192,  14'd1671,  -14'd367,  14'd366,  14'd325,  
-14'd87,  14'd472,  -14'd1636,  -14'd1073,  -14'd1446,  -14'd584,  -14'd319,  -14'd1881,  14'd956,  14'd1171,  14'd269,  14'd86,  14'd206,  14'd401,  -14'd1185,  14'd593,  
14'd1054,  14'd167,  -14'd1456,  -14'd297,  -14'd319,  -14'd398,  14'd563,  14'd1218,  
-14'd569,  14'd678,  -14'd884,  14'd724,  14'd682,  14'd970,  -14'd418,  -14'd1409,  14'd779,  14'd986,  14'd508,  14'd726,  14'd1259,  14'd887,  -14'd1007,  14'd280,  
-14'd131,  14'd762,  14'd725,  14'd1516,  -14'd132,  14'd1078,  -14'd781,  -14'd1672,  -14'd1153,  14'd1447,  -14'd1531,  14'd601,  -14'd385,  -14'd968,  -14'd220,  -14'd990,  
14'd427,  14'd1367,  -14'd1044,  14'd136,  14'd1576,  14'd896,  -14'd1433,  -14'd491,  -14'd982,  14'd1445,  -14'd1113,  14'd578,  -14'd445,  14'd800,  14'd294,  14'd103,  
14'd585,  -14'd761,  -14'd217,  14'd1134,  14'd44,  14'd1289,  -14'd33,  -14'd491,  -14'd110,  -14'd891,  -14'd1495,  -14'd333,  14'd554,  14'd411,  14'd2111,  -14'd423,  
-14'd524,  -14'd1154,  14'd228,  -14'd167,  14'd233,  14'd994,  14'd307,  14'd1723,  14'd127,  -14'd741,  -14'd1370,  -14'd1816,  -14'd1054,  -14'd807,  14'd531,  14'd1987,  
14'd120,  14'd858,  14'd28,  -14'd799,  14'd370,  14'd1409,  -14'd1731,  14'd1256,  14'd96,  -14'd1514,  14'd1490,  -14'd1338,  14'd1105,  -14'd665,  14'd674,  -14'd132,  
-14'd1084,  -14'd395,  -14'd491,  14'd673,  -14'd489,  14'd1580,  14'd977,  14'd1492,  -14'd423,  14'd279,  -14'd1018,  14'd371,  14'd348,  -14'd1910,  14'd779,  14'd1339,  
-14'd1627,  14'd1460,  14'd755,  14'd709,  -14'd54,  -14'd462,  14'd549,  14'd306,  
-14'd99,  14'd141,  -14'd2089,  14'd1421,  -14'd397,  -14'd1310,  14'd1371,  -14'd229,  14'd183,  -14'd112,  14'd1067,  14'd522,  14'd320,  14'd94,  -14'd396,  14'd1024,  
-14'd453,  14'd623,  14'd916,  14'd791,  -14'd398,  14'd759,  -14'd33,  14'd300,  14'd1502,  -14'd117,  14'd1691,  14'd753,  14'd179,  14'd629,  14'd560,  -14'd423,  
14'd969,  -14'd1,  -14'd984,  14'd1175,  -14'd1134,  14'd1922,  14'd843,  -14'd1223,  14'd914,  14'd304,  14'd385,  14'd699,  -14'd478,  14'd319,  14'd662,  14'd1713,  
-14'd295,  -14'd492,  14'd697,  -14'd770,  14'd1643,  -14'd112,  14'd1921,  14'd715,  14'd625,  14'd1353,  -14'd1339,  -14'd889,  -14'd506,  14'd1598,  14'd241,  -14'd991,  
-14'd373,  -14'd502,  -14'd494,  14'd1121,  14'd632,  -14'd104,  14'd242,  14'd467,  14'd617,  14'd1905,  -14'd526,  -14'd855,  -14'd23,  14'd209,  -14'd610,  14'd784,  
14'd1175,  14'd479,  -14'd1139,  14'd1589,  14'd419,  -14'd1186,  14'd182,  14'd1860,  14'd1449,  -14'd388,  -14'd197,  14'd823,  -14'd705,  -14'd556,  -14'd324,  -14'd420,  
14'd1225,  -14'd128,  -14'd796,  -14'd220,  -14'd432,  14'd31,  -14'd992,  14'd2043,  -14'd770,  14'd1071,  14'd514,  14'd567,  14'd880,  -14'd649,  14'd1458,  -14'd364,  
-14'd735,  14'd206,  -14'd186,  14'd706,  14'd1367,  -14'd292,  14'd872,  -14'd381,  
-14'd2408,  14'd507,  14'd878,  -14'd171,  -14'd2228,  14'd1042,  14'd201,  -14'd545,  -14'd1585,  -14'd1558,  14'd1150,  -14'd707,  -14'd1200,  14'd77,  14'd659,  14'd506,  
-14'd1461,  14'd255,  14'd355,  14'd341,  14'd674,  -14'd334,  14'd324,  -14'd1289,  -14'd650,  14'd76,  14'd1290,  14'd1076,  -14'd175,  14'd1000,  -14'd145,  -14'd853,  
-14'd925,  14'd136,  -14'd1060,  14'd66,  14'd2545,  14'd950,  -14'd1811,  14'd187,  14'd231,  14'd474,  14'd197,  -14'd81,  -14'd692,  14'd359,  14'd174,  14'd22,  
14'd414,  -14'd1066,  14'd1503,  -14'd1272,  14'd541,  14'd30,  -14'd479,  14'd104,  -14'd2508,  14'd884,  14'd1630,  -14'd573,  -14'd706,  -14'd485,  14'd1795,  14'd632,  
14'd1279,  14'd235,  14'd1237,  -14'd744,  -14'd123,  -14'd12,  14'd369,  14'd218,  14'd910,  -14'd2418,  14'd570,  14'd725,  -14'd28,  -14'd879,  -14'd326,  -14'd187,  
14'd67,  14'd976,  -14'd630,  -14'd1300,  14'd1411,  14'd1387,  14'd1218,  14'd617,  14'd806,  14'd45,  14'd917,  -14'd811,  -14'd8,  -14'd183,  14'd199,  14'd1612,  
14'd912,  14'd164,  14'd638,  -14'd1583,  14'd681,  -14'd1544,  14'd1201,  14'd393,  14'd274,  -14'd833,  -14'd421,  -14'd1010,  -14'd247,  14'd3698,  -14'd1278,  14'd449,  
-14'd937,  -14'd409,  -14'd207,  14'd97,  14'd221,  -14'd109,  -14'd1049,  14'd1588,  
-14'd2482,  14'd441,  -14'd547,  -14'd70,  14'd121,  14'd443,  14'd1423,  14'd54,  14'd2236,  14'd63,  14'd1832,  14'd322,  14'd1498,  14'd372,  -14'd617,  14'd129,  
-14'd1102,  -14'd22,  14'd1349,  14'd1519,  -14'd792,  14'd1630,  -14'd1049,  -14'd1348,  -14'd614,  -14'd375,  14'd200,  14'd1221,  -14'd252,  14'd100,  14'd711,  -14'd1321,  
-14'd886,  -14'd474,  -14'd407,  14'd1261,  -14'd692,  -14'd106,  14'd680,  -14'd138,  -14'd336,  14'd1014,  -14'd1387,  -14'd30,  -14'd858,  14'd219,  14'd778,  14'd2154,  
-14'd570,  14'd357,  14'd1393,  -14'd389,  -14'd730,  -14'd962,  -14'd415,  -14'd471,  -14'd675,  14'd340,  14'd189,  -14'd1170,  14'd939,  -14'd217,  14'd1256,  14'd222,  
-14'd787,  14'd143,  14'd369,  14'd1731,  14'd192,  14'd933,  14'd700,  14'd879,  14'd469,  -14'd1060,  14'd96,  14'd238,  -14'd1459,  14'd696,  -14'd1059,  14'd731,  
14'd839,  14'd473,  -14'd112,  14'd174,  14'd731,  14'd396,  14'd1197,  14'd356,  -14'd234,  14'd723,  14'd62,  14'd930,  -14'd282,  14'd256,  -14'd10,  -14'd352,  
14'd258,  14'd900,  -14'd188,  14'd161,  -14'd1577,  14'd438,  -14'd633,  14'd1656,  -14'd765,  14'd1308,  -14'd132,  -14'd747,  -14'd1150,  14'd2171,  -14'd339,  14'd164,  
-14'd242,  -14'd1015,  14'd1781,  14'd1327,  -14'd752,  14'd436,  -14'd647,  -14'd114,  
14'd935,  -14'd353,  14'd999,  14'd595,  14'd527,  -14'd875,  -14'd685,  -14'd614,  -14'd138,  14'd591,  -14'd210,  -14'd1692,  14'd1407,  14'd723,  14'd1314,  14'd0,  
-14'd178,  14'd369,  -14'd101,  -14'd576,  14'd1009,  -14'd42,  -14'd1027,  14'd533,  14'd452,  14'd91,  -14'd395,  -14'd956,  14'd1067,  14'd894,  14'd1265,  14'd1627,  
14'd141,  14'd227,  -14'd1011,  -14'd238,  14'd1260,  14'd440,  14'd1811,  -14'd1849,  -14'd722,  14'd1297,  -14'd417,  -14'd395,  -14'd552,  14'd121,  -14'd1482,  -14'd1044,  
-14'd298,  14'd825,  14'd187,  14'd37,  14'd1610,  14'd1004,  -14'd1540,  14'd757,  14'd406,  -14'd1316,  14'd332,  14'd520,  14'd608,  14'd162,  -14'd845,  -14'd996,  
14'd1477,  14'd158,  14'd258,  -14'd341,  -14'd612,  14'd1175,  14'd939,  -14'd249,  14'd105,  -14'd803,  14'd535,  -14'd1039,  14'd152,  14'd1037,  -14'd745,  -14'd26,  
14'd320,  -14'd316,  -14'd974,  14'd2285,  14'd1162,  -14'd33,  14'd329,  14'd346,  -14'd1641,  -14'd401,  -14'd27,  -14'd1767,  14'd505,  14'd803,  -14'd761,  -14'd1296,  
-14'd405,  14'd500,  -14'd1140,  -14'd85,  -14'd1140,  14'd812,  -14'd258,  14'd623,  -14'd1332,  14'd1237,  -14'd125,  14'd1437,  -14'd716,  -14'd302,  14'd1368,  14'd567,  
-14'd139,  -14'd219,  14'd375,  -14'd36,  -14'd28,  14'd268,  -14'd237,  -14'd41,  
-14'd1895,  -14'd1370,  14'd1858,  -14'd715,  -14'd851,  -14'd811,  -14'd142,  14'd1630,  14'd43,  14'd855,  14'd2764,  14'd18,  -14'd573,  14'd936,  -14'd1313,  14'd1211,  
-14'd1386,  14'd579,  14'd1182,  -14'd1104,  -14'd485,  -14'd198,  -14'd9,  14'd245,  14'd1130,  14'd711,  14'd590,  14'd652,  -14'd673,  -14'd345,  -14'd1238,  14'd342,  
14'd897,  14'd910,  -14'd388,  14'd726,  14'd178,  14'd1477,  -14'd675,  14'd1506,  -14'd129,  14'd1363,  14'd768,  14'd1126,  14'd1371,  14'd1104,  -14'd262,  14'd200,  
-14'd521,  14'd828,  14'd1062,  14'd635,  14'd170,  -14'd1738,  14'd429,  14'd1377,  14'd816,  -14'd1177,  14'd1173,  14'd922,  -14'd749,  -14'd336,  14'd749,  14'd1662,  
14'd221,  14'd752,  -14'd1,  -14'd119,  -14'd578,  -14'd502,  14'd694,  -14'd191,  -14'd5,  -14'd248,  14'd281,  -14'd617,  -14'd328,  -14'd1089,  14'd920,  -14'd347,  
-14'd861,  -14'd408,  14'd152,  -14'd938,  14'd725,  14'd34,  -14'd122,  14'd274,  14'd1259,  14'd371,  14'd1112,  14'd570,  -14'd1268,  14'd150,  -14'd378,  14'd824,  
14'd21,  14'd1727,  14'd492,  14'd603,  -14'd292,  -14'd128,  -14'd659,  14'd1452,  14'd867,  -14'd598,  -14'd832,  -14'd680,  14'd746,  14'd1830,  -14'd175,  -14'd569,  
14'd694,  -14'd1033,  -14'd619,  14'd188,  14'd442,  -14'd176,  -14'd331,  14'd1114,  
14'd759,  -14'd855,  -14'd358,  14'd91,  14'd532,  -14'd936,  -14'd801,  14'd836,  -14'd455,  14'd599,  -14'd2038,  14'd456,  14'd197,  -14'd29,  14'd1287,  -14'd1487,  
14'd257,  -14'd214,  -14'd2778,  -14'd428,  14'd1122,  -14'd341,  -14'd617,  -14'd1033,  -14'd1132,  14'd486,  14'd133,  -14'd1313,  -14'd456,  14'd1615,  14'd629,  -14'd176,  
14'd935,  14'd1427,  -14'd609,  14'd954,  14'd958,  14'd512,  -14'd1053,  -14'd1854,  14'd159,  14'd323,  14'd713,  -14'd2806,  14'd1465,  14'd111,  -14'd1130,  -14'd1155,  
-14'd1105,  -14'd476,  14'd1426,  -14'd1878,  -14'd1003,  14'd1575,  -14'd418,  14'd660,  -14'd1077,  -14'd64,  -14'd1786,  14'd862,  -14'd777,  -14'd1419,  14'd872,  14'd241,  
14'd152,  14'd555,  -14'd290,  -14'd919,  -14'd1236,  14'd69,  14'd770,  -14'd795,  -14'd800,  14'd577,  14'd325,  14'd417,  14'd145,  14'd1012,  14'd410,  14'd422,  
14'd532,  -14'd1755,  -14'd974,  -14'd277,  14'd724,  14'd60,  14'd150,  14'd583,  -14'd1986,  14'd402,  14'd481,  -14'd1687,  -14'd98,  14'd1333,  -14'd1292,  14'd712,  
-14'd440,  14'd645,  -14'd291,  -14'd1299,  14'd1529,  -14'd179,  -14'd377,  14'd631,  -14'd193,  -14'd405,  -14'd1011,  -14'd496,  -14'd862,  14'd20,  -14'd330,  14'd1774,  
-14'd1305,  14'd1002,  14'd310,  14'd531,  -14'd1000,  -14'd904,  14'd602,  -14'd201,  
14'd234,  -14'd818,  14'd1047,  -14'd34,  14'd338,  14'd120,  14'd718,  -14'd230,  14'd427,  -14'd881,  14'd241,  14'd411,  -14'd1444,  14'd222,  -14'd1104,  -14'd1079,  
14'd1135,  14'd877,  14'd1187,  14'd838,  -14'd784,  -14'd121,  14'd501,  -14'd166,  14'd1267,  14'd565,  -14'd791,  -14'd501,  -14'd132,  14'd1200,  -14'd1254,  -14'd1635,  
-14'd156,  14'd155,  14'd308,  14'd139,  -14'd945,  14'd1125,  14'd139,  14'd1399,  14'd532,  14'd300,  14'd920,  -14'd872,  -14'd828,  -14'd40,  14'd222,  14'd1409,  
14'd17,  14'd645,  -14'd925,  14'd779,  -14'd2011,  -14'd563,  14'd1681,  -14'd1066,  14'd472,  14'd827,  14'd51,  -14'd921,  14'd325,  -14'd1123,  -14'd32,  -14'd711,  
-14'd535,  14'd599,  14'd125,  -14'd550,  14'd629,  14'd792,  14'd145,  14'd504,  -14'd293,  14'd75,  14'd10,  -14'd1653,  14'd119,  14'd564,  -14'd130,  -14'd1394,  
-14'd545,  -14'd1071,  14'd1256,  14'd1769,  14'd1171,  14'd766,  -14'd378,  -14'd1173,  14'd1207,  14'd1253,  14'd954,  -14'd287,  -14'd1525,  14'd1812,  -14'd734,  14'd1207,  
-14'd577,  -14'd447,  14'd1075,  14'd998,  -14'd110,  14'd108,  14'd683,  14'd1807,  -14'd467,  14'd78,  -14'd388,  14'd626,  14'd434,  -14'd1682,  14'd1735,  -14'd1266,  
-14'd1411,  -14'd1026,  14'd205,  14'd278,  14'd733,  -14'd365,  -14'd299,  -14'd548,  
-14'd658,  14'd894,  -14'd1910,  14'd1105,  14'd443,  -14'd152,  -14'd124,  14'd162,  14'd231,  -14'd1083,  -14'd1735,  14'd967,  14'd1787,  -14'd1021,  -14'd693,  14'd4,  
-14'd177,  14'd64,  -14'd166,  -14'd85,  -14'd171,  14'd117,  14'd90,  -14'd220,  -14'd349,  -14'd1660,  14'd830,  14'd230,  14'd239,  -14'd608,  14'd1329,  -14'd1510,  
-14'd426,  -14'd728,  -14'd377,  14'd660,  -14'd1497,  14'd359,  14'd1386,  -14'd294,  14'd843,  -14'd573,  -14'd1318,  14'd296,  14'd476,  -14'd847,  14'd529,  14'd1546,  
-14'd981,  -14'd2292,  -14'd289,  -14'd666,  14'd1029,  14'd1090,  -14'd1591,  -14'd183,  14'd1147,  14'd462,  -14'd488,  -14'd1559,  14'd2020,  -14'd308,  14'd386,  -14'd336,  
14'd50,  14'd130,  -14'd769,  -14'd335,  14'd1478,  -14'd467,  14'd494,  14'd1559,  -14'd777,  14'd991,  -14'd305,  14'd1559,  14'd782,  14'd1445,  -14'd1192,  -14'd364,  
14'd816,  14'd1258,  -14'd1537,  14'd728,  -14'd1238,  14'd58,  14'd768,  14'd1413,  14'd353,  14'd69,  14'd95,  14'd376,  -14'd371,  -14'd1,  -14'd722,  14'd1665,  
-14'd344,  14'd145,  14'd933,  14'd1327,  14'd174,  -14'd569,  14'd1209,  14'd1615,  -14'd630,  -14'd256,  14'd457,  14'd1971,  14'd304,  -14'd68,  14'd885,  14'd566,  
-14'd152,  14'd1763,  14'd1031,  14'd208,  14'd1539,  -14'd1276,  14'd194,  -14'd296
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule


module bias_fc3_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC3-1][0:`OUTPUT_NUM_FC3-1][`WD_BIAS:0] weight	 = {
-24'd186531,  24'd166143,  -24'd211411,  -24'd80228,  -24'd155665,  24'd207658,  -24'd315652,  -24'd209780,  24'd326774,  24'd153726
	};

	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule




module wieght_fc3_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3*`OUTPUT_BATCH_FC3)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC2*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC3*`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3-1][0:`OUTPUT_NUM_FC3-1][0:`OUTPUT_NUM_FC2-1][`WD:0] weight	 = {
-14'd98,  14'd854,  -14'd128,  -14'd253,  14'd282,  14'd458,  14'd239,  -14'd218,  -14'd929,  -14'd722,  14'd2043,  -14'd1381,  -14'd454,  -14'd79,  -14'd1025,  14'd817,  
14'd1185,  14'd191,  -14'd193,  14'd2087,  14'd2594,  -14'd1959,  -14'd1373,  -14'd177,  -14'd1614,  14'd1310,  14'd501,  -14'd154,  -14'd745,  14'd999,  14'd341,  14'd1235,  
-14'd1175,  -14'd1978,  -14'd687,  -14'd1884,  -14'd526,  14'd703,  14'd505,  -14'd517,  14'd773,  -14'd142,  14'd1461,  -14'd682,  -14'd1755,  14'd352,  -14'd366,  14'd328,  
-14'd2046,  -14'd266,  14'd1195,  14'd323,  14'd2046,  -14'd725,  -14'd1261,  14'd1157,  -14'd753,  14'd2069,  14'd4,  -14'd260,  -14'd468,  -14'd482,  14'd366,  -14'd1159,  
14'd1714,  -14'd1828,  -14'd485,  -14'd350,  -14'd929,  -14'd1023,  -14'd77,  -14'd2441,  -14'd112,  -14'd547,  -14'd931,  14'd301,  14'd195,  -14'd712,  14'd1202,  -14'd392,  
-14'd472,  -14'd1170,  14'd1552,  -14'd1047,  
14'd1141,  -14'd1711,  14'd333,  -14'd793,  -14'd115,  14'd423,  14'd858,  -14'd648,  -14'd146,  -14'd1044,  -14'd1922,  14'd958,  14'd118,  14'd1378,  14'd506,  14'd499,  
-14'd1158,  14'd1050,  -14'd1035,  -14'd795,  14'd1780,  -14'd549,  -14'd52,  14'd142,  -14'd1750,  -14'd201,  -14'd339,  14'd1316,  14'd994,  -14'd204,  14'd1351,  -14'd454,  
14'd19,  -14'd1073,  -14'd8,  14'd1609,  -14'd900,  -14'd987,  -14'd510,  -14'd1577,  14'd1217,  -14'd775,  -14'd2298,  -14'd1737,  14'd1120,  14'd784,  -14'd7,  14'd784,  
-14'd855,  14'd1387,  -14'd1959,  -14'd864,  -14'd273,  14'd803,  14'd2088,  -14'd989,  -14'd523,  -14'd632,  -14'd2315,  14'd2014,  -14'd1021,  14'd240,  -14'd1424,  -14'd452,  
14'd1572,  -14'd945,  14'd512,  14'd2238,  14'd736,  -14'd1466,  -14'd1002,  14'd1244,  14'd931,  14'd260,  -14'd1607,  -14'd901,  -14'd95,  -14'd1688,  -14'd1404,  14'd513,  
14'd850,  -14'd2014,  14'd2011,  -14'd315,  
-14'd1414,  -14'd1437,  14'd916,  -14'd194,  14'd1932,  14'd790,  -14'd792,  14'd191,  14'd540,  -14'd769,  14'd935,  14'd1696,  14'd315,  -14'd1332,  -14'd488,  -14'd637,  
-14'd276,  -14'd2523,  -14'd1319,  14'd836,  14'd1597,  14'd217,  -14'd649,  -14'd1355,  14'd106,  -14'd429,  -14'd175,  -14'd493,  -14'd772,  14'd1492,  -14'd2653,  -14'd111,  
-14'd2471,  -14'd487,  14'd107,  -14'd1318,  14'd340,  14'd1153,  14'd392,  14'd1810,  -14'd108,  -14'd379,  14'd376,  -14'd817,  14'd113,  -14'd203,  14'd924,  14'd823,  
14'd1050,  14'd1196,  -14'd2247,  -14'd1737,  -14'd515,  -14'd594,  -14'd849,  -14'd685,  14'd335,  14'd1207,  14'd31,  14'd426,  -14'd143,  -14'd1687,  -14'd126,  14'd1280,  
14'd587,  -14'd1306,  14'd419,  -14'd970,  -14'd560,  14'd633,  14'd598,  14'd355,  -14'd1146,  14'd705,  -14'd940,  14'd164,  -14'd376,  14'd1700,  14'd433,  -14'd1289,  
14'd1893,  -14'd404,  -14'd107,  -14'd972,  
-14'd10,  -14'd893,  14'd132,  -14'd1917,  14'd1106,  14'd169,  -14'd987,  -14'd847,  14'd345,  -14'd600,  -14'd1285,  -14'd1000,  14'd1903,  -14'd1144,  -14'd1134,  14'd359,  
-14'd1117,  14'd566,  -14'd764,  14'd1514,  -14'd2527,  -14'd1013,  -14'd1114,  -14'd1500,  -14'd119,  14'd408,  -14'd1206,  14'd377,  -14'd1323,  14'd961,  -14'd260,  -14'd376,  
14'd136,  14'd510,  -14'd1088,  14'd1011,  14'd583,  -14'd899,  -14'd349,  14'd993,  -14'd862,  -14'd441,  14'd1333,  14'd647,  14'd1128,  -14'd1577,  -14'd592,  -14'd971,  
14'd1208,  -14'd1891,  14'd203,  14'd1395,  -14'd1323,  -14'd38,  -14'd471,  -14'd766,  -14'd808,  -14'd696,  14'd916,  14'd67,  14'd176,  14'd286,  -14'd153,  14'd457,  
-14'd1533,  14'd2594,  -14'd260,  14'd687,  14'd45,  14'd43,  -14'd1587,  14'd1229,  -14'd1860,  14'd821,  -14'd568,  14'd18,  14'd1153,  14'd124,  14'd9,  -14'd477,  
-14'd1772,  -14'd466,  14'd282,  14'd2047,  
-14'd1185,  14'd1312,  14'd62,  14'd453,  -14'd1288,  14'd775,  14'd2078,  14'd1111,  -14'd1625,  -14'd17,  -14'd581,  -14'd987,  -14'd663,  14'd1471,  14'd832,  -14'd1494,  
14'd1432,  -14'd826,  -14'd1952,  -14'd298,  -14'd1327,  14'd696,  -14'd201,  -14'd2033,  14'd846,  -14'd413,  -14'd3036,  -14'd472,  14'd1688,  14'd624,  -14'd1579,  -14'd1267,  
14'd30,  -14'd1673,  -14'd400,  14'd147,  -14'd1340,  14'd885,  14'd1068,  -14'd1773,  14'd11,  -14'd512,  14'd107,  14'd1708,  14'd416,  14'd1023,  -14'd296,  14'd372,  
14'd796,  -14'd533,  14'd887,  -14'd840,  14'd982,  14'd9,  -14'd705,  -14'd344,  -14'd242,  14'd382,  -14'd709,  14'd1604,  -14'd77,  -14'd291,  -14'd1244,  14'd1176,  
14'd418,  -14'd1606,  14'd156,  14'd1588,  -14'd1963,  -14'd965,  14'd1359,  -14'd905,  -14'd1781,  -14'd1427,  14'd960,  14'd1401,  -14'd1642,  14'd924,  -14'd1694,  14'd1284,  
-14'd1282,  14'd928,  -14'd1079,  -14'd1271,  
14'd2227,  14'd1116,  -14'd1479,  -14'd1476,  14'd2026,  -14'd1255,  -14'd1537,  14'd504,  14'd1177,  14'd1207,  14'd460,  14'd2044,  -14'd1391,  -14'd1186,  14'd178,  -14'd720,  
14'd591,  14'd1505,  14'd853,  14'd827,  -14'd1231,  14'd641,  -14'd925,  14'd1346,  14'd1255,  14'd696,  14'd901,  14'd200,  -14'd684,  14'd57,  14'd450,  -14'd640,  
-14'd26,  -14'd236,  14'd570,  14'd2151,  -14'd1220,  -14'd2257,  -14'd1820,  14'd519,  14'd816,  14'd65,  -14'd1355,  -14'd1122,  -14'd1331,  -14'd893,  -14'd632,  14'd0,  
14'd1237,  14'd1354,  14'd175,  14'd1232,  14'd477,  -14'd1810,  -14'd2056,  14'd514,  -14'd691,  -14'd434,  14'd544,  -14'd1398,  14'd7,  14'd55,  14'd92,  -14'd1535,  
-14'd91,  -14'd360,  14'd1365,  14'd357,  -14'd175,  -14'd901,  -14'd664,  -14'd142,  14'd2039,  -14'd169,  14'd1137,  14'd518,  14'd508,  -14'd387,  14'd48,  14'd1085,  
-14'd1500,  14'd675,  -14'd1436,  14'd324,  
14'd1854,  -14'd1011,  -14'd224,  -14'd59,  -14'd95,  -14'd1304,  -14'd229,  14'd1097,  14'd412,  14'd1112,  -14'd785,  -14'd1125,  -14'd3030,  -14'd175,  -14'd1220,  -14'd1174,  
14'd1142,  -14'd437,  -14'd1523,  -14'd1041,  14'd334,  14'd353,  -14'd1449,  -14'd715,  14'd754,  -14'd613,  -14'd56,  14'd42,  -14'd1697,  14'd199,  14'd1110,  14'd710,  
-14'd692,  14'd1741,  -14'd126,  -14'd523,  -14'd1485,  -14'd1280,  14'd807,  -14'd818,  -14'd636,  -14'd1471,  14'd2170,  -14'd1810,  14'd150,  -14'd558,  14'd787,  -14'd121,  
-14'd518,  -14'd1566,  14'd1064,  -14'd958,  14'd98,  14'd905,  14'd268,  14'd771,  -14'd3,  14'd401,  14'd627,  -14'd25,  14'd647,  -14'd1435,  14'd657,  -14'd1864,  
14'd557,  14'd924,  -14'd258,  14'd101,  -14'd106,  14'd415,  14'd638,  -14'd1033,  14'd979,  -14'd704,  14'd444,  -14'd1423,  -14'd1081,  14'd649,  -14'd1001,  14'd251,  
14'd528,  14'd807,  -14'd812,  -14'd2450,  
-14'd1413,  -14'd326,  14'd689,  -14'd2698,  -14'd1103,  14'd700,  -14'd2262,  -14'd688,  -14'd878,  -14'd759,  -14'd2256,  14'd448,  14'd339,  14'd629,  -14'd957,  14'd133,  
14'd901,  -14'd90,  -14'd928,  -14'd604,  -14'd532,  -14'd680,  -14'd853,  -14'd797,  -14'd429,  -14'd178,  -14'd214,  -14'd757,  14'd1814,  -14'd394,  14'd606,  -14'd91,  
14'd42,  -14'd354,  14'd2232,  -14'd713,  14'd256,  14'd1676,  -14'd1353,  -14'd502,  -14'd558,  14'd330,  -14'd2260,  -14'd63,  14'd1630,  14'd1660,  -14'd678,  -14'd314,  
14'd245,  14'd440,  14'd667,  -14'd1540,  14'd761,  14'd267,  14'd148,  -14'd1128,  14'd627,  -14'd2627,  -14'd1530,  14'd962,  -14'd196,  14'd1344,  -14'd1010,  -14'd980,  
-14'd235,  14'd2088,  14'd62,  -14'd2374,  14'd1464,  -14'd649,  14'd187,  14'd73,  14'd235,  -14'd235,  14'd650,  14'd273,  14'd1034,  14'd824,  14'd1068,  -14'd83,  
14'd699,  -14'd1524,  14'd349,  14'd8,  
14'd102,  14'd1049,  14'd774,  -14'd222,  -14'd37,  -14'd58,  14'd13,  -14'd834,  -14'd273,  14'd2089,  -14'd1694,  -14'd2010,  14'd243,  -14'd1573,  -14'd83,  14'd269,  
14'd471,  14'd616,  14'd978,  14'd258,  14'd139,  14'd1182,  -14'd199,  -14'd760,  14'd120,  -14'd930,  -14'd1502,  14'd169,  -14'd1136,  -14'd801,  -14'd2220,  -14'd962,  
-14'd1468,  14'd927,  -14'd809,  14'd892,  14'd259,  14'd151,  -14'd245,  14'd573,  -14'd153,  14'd247,  -14'd1019,  14'd1882,  -14'd1408,  14'd1301,  14'd251,  14'd287,  
-14'd1344,  -14'd1893,  -14'd1276,  14'd1161,  14'd1059,  14'd1041,  14'd645,  14'd520,  -14'd288,  -14'd1213,  14'd339,  -14'd1269,  14'd1391,  -14'd1259,  14'd1138,  -14'd2,  
14'd955,  14'd1208,  -14'd1243,  -14'd769,  14'd52,  -14'd1768,  -14'd1563,  14'd16,  14'd843,  14'd95,  14'd543,  -14'd1853,  -14'd1253,  14'd159,  14'd339,  -14'd1919,  
14'd1265,  14'd1797,  -14'd59,  -14'd350,  
14'd393,  14'd505,  14'd746,  14'd401,  14'd710,  -14'd864,  14'd674,  14'd591,  -14'd786,  -14'd1103,  14'd651,  14'd830,  14'd1246,  14'd1391,  14'd808,  14'd426,  
-14'd1605,  -14'd133,  -14'd450,  -14'd708,  -14'd21,  -14'd758,  14'd1077,  14'd266,  14'd1183,  -14'd404,  14'd437,  -14'd587,  14'd589,  -14'd2290,  -14'd1123,  -14'd481,  
14'd206,  -14'd1457,  14'd405,  -14'd176,  -14'd820,  14'd1635,  14'd604,  14'd1264,  14'd1414,  14'd1276,  -14'd574,  14'd271,  14'd739,  -14'd248,  14'd297,  -14'd138,  
-14'd2288,  -14'd733,  -14'd192,  14'd816,  14'd884,  -14'd164,  -14'd2642,  -14'd133,  -14'd265,  14'd1110,  14'd680,  -14'd1942,  14'd190,  14'd946,  14'd2297,  14'd1141,  
-14'd482,  -14'd2955,  14'd543,  14'd246,  -14'd24,  14'd1551,  14'd1316,  14'd1020,  -14'd569,  -14'd2639,  14'd1300,  -14'd1677,  -14'd243,  -14'd1848,  -14'd1329,  14'd442,  
-14'd1629,  -14'd1329,  -14'd570,  -14'd45
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule

