// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION
`include "global.v"


module bias_conv1_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV1-1][0:`OUTPUT_NUM_CONV1-1][`WD_BIAS:0] weight	 = {	
		-24'd33091,  -24'd345382,  -24'd986031,  -24'd314271,  24'd400309,  -24'd448129
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_conv1_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV1*`KERNEL_SIZE_CONV1-1][0:`OUTPUT_NUM_CONV1-1][12:0] weight	 = {
13'd123,  13'd232,  -13'd455,  13'd444,  -13'd794,  -13'd1534,  
13'd475,  -13'd381,  -13'd258,  -13'd171,  -13'd986,  -13'd940,  
-13'd973,  -13'd682,  -13'd184,  13'd257,  -13'd1381,  13'd35,  
-13'd958,  -13'd187,  13'd457,  13'd532,  -13'd1075,  13'd428,  
-13'd1568,  13'd505,  13'd123,  -13'd333,  -13'd1129,  13'd1181,  

13'd844,  -13'd388,  -13'd645,  13'd1049,  -13'd89,  -13'd1103,  
13'd104,  -13'd577,  -13'd209,  13'd512,  -13'd1471,  13'd355,  
13'd462,  13'd50,  13'd508,  13'd699,  -13'd887,  13'd650,  
-13'd621,  13'd481,  13'd790,  13'd952,  -13'd498,  13'd1062,  
-13'd1395,  13'd1,  13'd311,  -13'd665,  -13'd904,  -13'd335,  

13'd443,  -13'd192,  -13'd847,  13'd859,  13'd177,  -13'd416,  
13'd1275,  13'd106,  13'd493,  13'd444,  13'd372,  13'd355,  
13'd1281,  -13'd128,  13'd714,  13'd676,  13'd208,  13'd1024,  
13'd388,  13'd877,  13'd979,  13'd749,  13'd249,  13'd489,  
13'd626,  13'd559,  -13'd291,  13'd159,  13'd957,  -13'd1036,  

-13'd867,  -13'd189,  -13'd103,  -13'd3,  13'd1323,  13'd81,  
13'd734,  13'd175,  13'd262,  13'd652,  13'd1271,  13'd519,  
13'd37,  13'd1121,  13'd1490,  13'd839,  13'd967,  13'd884,  
13'd1062,  13'd1010,  13'd84,  13'd1205,  13'd1151,  -13'd54,  
13'd360,  -13'd295,  -13'd700,  13'd1154,  13'd622,  -13'd1790,  

-13'd762,  13'd41,  13'd931,  13'd3,  13'd853,  13'd221,  
-13'd530,  13'd554,  13'd722,  -13'd890,  13'd232,  13'd16,  
-13'd367,  13'd26,  13'd667,  -13'd9,  13'd689,  13'd613,  
13'd574,  13'd1025,  -13'd416,  13'd200,  -13'd111,  -13'd108,  
-13'd221,  13'd731,  -13'd629,  13'd985,  13'd217,  -13'd941
		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule	


module bias_conv2_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV2-1][0:`OUTPUT_NUM_CONV2-1][`WD_BIAS:0] weight	 = {
	-24'd492928,  -24'd252352,  24'd425549,  -24'd126681,  -24'd362367,  -24'd84127,  24'd122339,  -24'd193094,  24'd178645,  24'd56283,  -24'd15047,  -24'd647019,  -24'd375850,  24'd168062,  -24'd242871,  -24'd1026233		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule



module wieght_conv2_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][`WD:0] weight	 = {
13'd467,  -13'd260,  13'd530,  13'd252,  -13'd156,  13'd527,  
-13'd711,  -13'd534,  13'd407,  13'd228,  -13'd443,  -13'd539,  
13'd638,  -13'd704,  -13'd978,  -13'd525,  -13'd6,  13'd214,  
-13'd29,  13'd201,  -13'd738,  -13'd249,  -13'd409,  -13'd1115,  
13'd236,  -13'd680,  -13'd226,  -13'd697,  -13'd622,  13'd122,  
-13'd726,  -13'd415,  13'd281,  -13'd111,  -13'd397,  13'd428,  
13'd136,  13'd174,  -13'd411,  13'd500,  -13'd318,  13'd126,  
13'd63,  13'd28,  -13'd620,  13'd135,  -13'd696,  13'd149,  
13'd122,  -13'd1082,  -13'd622,  -13'd306,  13'd387,  -13'd492,  
13'd740,  -13'd986,  -13'd982,  -13'd13,  -13'd1427,  13'd548,  
-13'd535,  -13'd320,  -13'd38,  -13'd151,  -13'd60,  -13'd1093,  
-13'd358,  -13'd293,  -13'd645,  -13'd3,  13'd229,  13'd184,  
-13'd217,  -13'd446,  -13'd219,  -13'd246,  13'd112,  13'd413,  
13'd600,  13'd131,  -13'd314,  13'd929,  13'd63,  -13'd140,  
13'd60,  13'd459,  -13'd289,  13'd282,  13'd601,  -13'd667,  
-13'd342,  13'd242,  -13'd157,  -13'd148,  -13'd357,  -13'd19,  

-13'd280,  13'd22,  -13'd507,  -13'd763,  -13'd228,  -13'd319,  
13'd273,  -13'd281,  -13'd309,  13'd707,  -13'd429,  -13'd465,  
-13'd1343,  -13'd738,  -13'd24,  -13'd759,  -13'd384,  -13'd255,  
13'd171,  13'd57,  -13'd295,  -13'd562,  -13'd62,  13'd267,  
-13'd1033,  -13'd125,  13'd445,  -13'd183,  -13'd573,  13'd414,  
-13'd162,  13'd542,  -13'd267,  13'd73,  -13'd146,  -13'd724,  
-13'd580,  13'd548,  -13'd231,  13'd707,  -13'd102,  13'd595,  
-13'd284,  -13'd295,  -13'd516,  13'd343,  -13'd25,  13'd121,  
-13'd272,  -13'd194,  13'd152,  -13'd545,  13'd32,  -13'd518,  
-13'd40,  -13'd1012,  13'd604,  -13'd28,  -13'd990,  13'd154,  
-13'd225,  -13'd411,  13'd271,  -13'd270,  13'd877,  13'd58,  
-13'd881,  -13'd11,  -13'd738,  13'd344,  13'd255,  -13'd35,  
13'd511,  -13'd92,  13'd242,  -13'd784,  -13'd113,  -13'd714,  
-13'd66,  -13'd816,  13'd632,  -13'd52,  13'd650,  -13'd57,  
13'd331,  13'd194,  13'd694,  -13'd31,  13'd233,  -13'd659,  
-13'd291,  13'd488,  -13'd153,  -13'd126,  13'd42,  -13'd462,  

-13'd17,  -13'd233,  13'd92,  -13'd745,  -13'd134,  -13'd595,  
13'd670,  -13'd598,  -13'd495,  13'd237,  -13'd161,  13'd100,  
-13'd519,  -13'd231,  -13'd604,  13'd799,  -13'd887,  -13'd601,  
13'd316,  -13'd115,  13'd283,  -13'd415,  -13'd25,  13'd711,  
-13'd269,  -13'd417,  13'd117,  13'd87,  -13'd1433,  -13'd263,  
13'd615,  13'd316,  13'd54,  13'd177,  -13'd158,  -13'd899,  
13'd148,  -13'd578,  -13'd29,  -13'd551,  13'd597,  13'd244,  
-13'd380,  13'd482,  13'd605,  13'd154,  -13'd581,  13'd350,  
-13'd582,  -13'd104,  -13'd607,  -13'd393,  -13'd507,  -13'd582,  
-13'd143,  -13'd807,  -13'd475,  -13'd368,  -13'd1232,  13'd406,  
13'd288,  13'd169,  -13'd346,  -13'd320,  13'd479,  -13'd920,  
13'd622,  -13'd491,  -13'd521,  13'd319,  13'd798,  -13'd438,  
-13'd629,  -13'd144,  -13'd550,  -13'd297,  -13'd10,  -13'd103,  
-13'd262,  -13'd235,  -13'd311,  -13'd300,  -13'd579,  -13'd616,  
-13'd59,  13'd576,  -13'd283,  13'd146,  13'd1198,  -13'd392,  
-13'd2,  13'd170,  -13'd30,  13'd572,  13'd357,  -13'd1455,  

13'd1201,  -13'd496,  -13'd690,  -13'd152,  -13'd452,  -13'd989,  
13'd225,  13'd676,  -13'd397,  13'd459,  -13'd296,  -13'd345,  
13'd331,  13'd147,  13'd480,  13'd197,  -13'd978,  13'd290,  
-13'd707,  -13'd821,  -13'd307,  -13'd837,  -13'd406,  13'd643,  
13'd439,  13'd78,  -13'd494,  13'd331,  -13'd1276,  -13'd1030,  
13'd253,  -13'd215,  -13'd149,  -13'd444,  13'd683,  -13'd835,  
-13'd373,  -13'd100,  -13'd186,  13'd256,  13'd312,  13'd515,  
13'd63,  -13'd298,  -13'd234,  13'd27,  -13'd215,  13'd657,  
-13'd19,  -13'd10,  -13'd69,  -13'd1017,  13'd506,  13'd346,  
-13'd183,  -13'd194,  13'd578,  -13'd599,  -13'd1210,  -13'd195,  
-13'd228,  13'd230,  13'd598,  -13'd78,  13'd317,  13'd135,  
13'd183,  -13'd429,  -13'd531,  13'd699,  -13'd175,  -13'd1257,  
-13'd538,  13'd147,  13'd313,  -13'd427,  -13'd23,  13'd32,  
-13'd979,  -13'd34,  -13'd228,  -13'd393,  -13'd1083,  -13'd577,  
-13'd125,  -13'd681,  -13'd209,  -13'd443,  13'd382,  -13'd476,  
13'd290,  13'd762,  -13'd435,  -13'd240,  13'd911,  -13'd333,  

13'd674,  -13'd26,  13'd334,  -13'd28,  13'd35,  13'd532,  
13'd709,  13'd104,  13'd52,  -13'd340,  13'd946,  -13'd27,  
-13'd86,  -13'd523,  13'd216,  13'd183,  -13'd374,  13'd460,  
-13'd391,  -13'd119,  13'd179,  -13'd500,  13'd42,  13'd596,  
13'd1078,  13'd336,  -13'd270,  13'd1333,  13'd851,  13'd164,  
-13'd226,  -13'd478,  -13'd305,  -13'd1509,  -13'd300,  13'd539,  
-13'd728,  -13'd615,  -13'd331,  13'd537,  -13'd223,  13'd1146,  
13'd138,  -13'd76,  -13'd426,  13'd116,  -13'd514,  -13'd77,  
-13'd308,  13'd467,  -13'd130,  -13'd426,  13'd279,  -13'd195,  
-13'd663,  13'd533,  13'd463,  13'd681,  -13'd429,  -13'd471,  
-13'd443,  13'd205,  13'd324,  13'd220,  -13'd440,  -13'd144,  
13'd715,  -13'd588,  -13'd981,  -13'd795,  13'd292,  -13'd1420,  
-13'd93,  13'd366,  13'd479,  13'd386,  -13'd448,  -13'd208,  
13'd665,  13'd619,  13'd867,  -13'd305,  -13'd912,  13'd974,  
-13'd198,  -13'd519,  13'd30,  -13'd357,  13'd696,  13'd63,  
-13'd152,  13'd189,  13'd165,  13'd38,  13'd668,  -13'd360,  


-13'd344,  13'd19,  13'd14,  -13'd680,  13'd20,  -13'd185,  
-13'd45,  -13'd426,  -13'd711,  -13'd801,  -13'd964,  -13'd720,  
13'd245,  -13'd298,  -13'd1,  -13'd481,  13'd639,  13'd128,  
-13'd423,  -13'd162,  -13'd676,  13'd174,  13'd137,  -13'd72,  
13'd538,  13'd48,  13'd217,  13'd212,  13'd414,  13'd740,  
-13'd219,  -13'd214,  -13'd492,  -13'd372,  -13'd149,  -13'd181,  
13'd112,  13'd21,  -13'd393,  -13'd169,  -13'd119,  -13'd306,  
13'd630,  13'd777,  -13'd327,  13'd432,  -13'd514,  -13'd565,  
-13'd329,  13'd45,  -13'd650,  -13'd578,  13'd186,  -13'd1304,  
-13'd543,  -13'd418,  -13'd784,  -13'd1046,  -13'd431,  13'd13,  
13'd41,  13'd697,  -13'd448,  13'd493,  13'd267,  -13'd496,  
-13'd239,  -13'd831,  -13'd214,  -13'd806,  13'd224,  13'd797,  
-13'd7,  13'd104,  -13'd152,  -13'd567,  -13'd524,  -13'd21,  
-13'd207,  13'd286,  13'd861,  13'd326,  13'd119,  13'd525,  
-13'd427,  -13'd453,  -13'd329,  13'd31,  -13'd576,  -13'd90,  
-13'd121,  -13'd518,  13'd574,  13'd262,  13'd497,  13'd315,  

13'd105,  13'd114,  -13'd382,  -13'd410,  -13'd671,  -13'd843,  
-13'd162,  13'd356,  13'd304,  13'd252,  -13'd682,  -13'd289,  
-13'd483,  -13'd428,  -13'd936,  -13'd188,  13'd60,  -13'd1326,  
13'd234,  13'd267,  13'd391,  13'd374,  -13'd182,  13'd208,  
13'd349,  -13'd350,  13'd739,  -13'd216,  13'd453,  13'd379,  
13'd356,  -13'd138,  13'd50,  13'd547,  -13'd740,  13'd188,  
-13'd64,  13'd185,  13'd982,  13'd159,  -13'd385,  -13'd95,  
13'd78,  -13'd531,  13'd200,  13'd374,  -13'd738,  -13'd330,  
13'd451,  13'd352,  13'd55,  -13'd514,  13'd103,  13'd353,  
-13'd247,  -13'd185,  -13'd898,  -13'd344,  -13'd500,  -13'd1461,  
13'd247,  13'd23,  13'd45,  13'd227,  13'd313,  -13'd596,  
13'd136,  -13'd44,  13'd192,  -13'd20,  -13'd154,  13'd523,  
-13'd307,  13'd605,  13'd620,  13'd81,  13'd24,  13'd450,  
13'd41,  -13'd271,  13'd481,  -13'd590,  13'd139,  13'd491,  
-13'd398,  13'd117,  13'd42,  13'd73,  -13'd229,  -13'd330,  
13'd701,  13'd677,  13'd203,  13'd52,  13'd944,  -13'd645,  

13'd284,  13'd909,  -13'd327,  13'd241,  -13'd220,  -13'd1063,  
13'd404,  -13'd77,  13'd112,  13'd277,  -13'd739,  -13'd121,  
-13'd643,  13'd508,  -13'd1,  13'd44,  -13'd947,  -13'd713,  
13'd691,  13'd108,  -13'd22,  13'd516,  -13'd299,  -13'd225,  
-13'd133,  13'd42,  13'd165,  -13'd835,  13'd616,  13'd695,  
13'd530,  13'd64,  13'd557,  13'd97,  13'd174,  -13'd753,  
13'd69,  13'd93,  13'd277,  -13'd48,  13'd14,  13'd462,  
13'd70,  -13'd119,  13'd803,  13'd267,  -13'd1508,  13'd6,  
-13'd111,  13'd133,  13'd429,  -13'd11,  13'd772,  13'd498,  
-13'd709,  13'd143,  -13'd284,  -13'd89,  13'd852,  13'd720,  
13'd467,  13'd84,  13'd95,  13'd580,  13'd518,  -13'd496,  
13'd254,  13'd428,  -13'd689,  -13'd505,  13'd622,  13'd498,  
-13'd618,  13'd490,  -13'd63,  13'd416,  13'd314,  13'd212,  
-13'd294,  -13'd469,  -13'd649,  -13'd531,  -13'd406,  -13'd398,  
-13'd79,  13'd664,  -13'd183,  13'd501,  -13'd642,  13'd87,  
13'd729,  13'd247,  13'd519,  13'd618,  13'd1363,  -13'd362,  

-13'd32,  -13'd131,  13'd772,  -13'd111,  -13'd310,  13'd401,  
13'd1018,  13'd406,  13'd170,  13'd330,  -13'd506,  13'd882,  
13'd840,  13'd1015,  13'd70,  13'd74,  -13'd403,  13'd977,  
13'd102,  13'd716,  13'd74,  13'd207,  -13'd404,  13'd646,  
-13'd261,  -13'd500,  13'd231,  -13'd446,  -13'd27,  13'd358,  
13'd604,  -13'd162,  -13'd501,  13'd525,  13'd63,  -13'd177,  
-13'd177,  13'd110,  13'd573,  -13'd455,  -13'd742,  13'd509,  
13'd65,  -13'd492,  13'd275,  13'd440,  -13'd821,  13'd465,  
-13'd316,  13'd651,  -13'd467,  13'd363,  13'd442,  -13'd816,  
-13'd370,  13'd610,  13'd511,  13'd52,  -13'd292,  13'd669,  
13'd785,  13'd321,  13'd363,  13'd94,  13'd1215,  -13'd41,  
13'd28,  13'd219,  -13'd140,  13'd358,  -13'd181,  -13'd547,  
13'd334,  -13'd393,  13'd483,  -13'd595,  -13'd33,  -13'd205,  
13'd220,  -13'd22,  13'd144,  -13'd477,  -13'd976,  13'd20,  
-13'd31,  -13'd180,  -13'd87,  13'd33,  -13'd598,  -13'd98,  
-13'd192,  13'd324,  -13'd279,  13'd707,  13'd640,  13'd47,  

13'd245,  -13'd504,  13'd970,  13'd636,  -13'd569,  13'd814,  
13'd357,  -13'd512,  13'd116,  -13'd60,  13'd309,  13'd500,  
13'd454,  -13'd846,  13'd77,  13'd276,  -13'd737,  13'd592,  
-13'd72,  -13'd363,  13'd164,  13'd189,  -13'd166,  13'd468,  
13'd223,  -13'd426,  -13'd551,  13'd532,  -13'd1446,  -13'd959,  
13'd28,  -13'd109,  13'd486,  13'd70,  -13'd308,  13'd608,  
-13'd435,  -13'd432,  -13'd489,  -13'd404,  -13'd1444,  13'd152,  
13'd74,  13'd592,  13'd326,  13'd137,  -13'd76,  -13'd165,  
-13'd256,  -13'd138,  13'd353,  13'd74,  13'd639,  13'd77,  
-13'd168,  -13'd211,  13'd396,  13'd443,  13'd100,  13'd647,  
13'd228,  13'd860,  13'd897,  -13'd406,  13'd650,  13'd726,  
13'd691,  -13'd662,  13'd8,  -13'd11,  -13'd818,  -13'd115,  
-13'd263,  -13'd324,  -13'd37,  13'd403,  13'd69,  13'd390,  
13'd374,  13'd124,  13'd175,  13'd419,  -13'd1306,  13'd447,  
13'd35,  13'd371,  13'd194,  13'd193,  13'd183,  13'd181,  
13'd307,  -13'd1163,  -13'd183,  13'd307,  -13'd34,  -13'd657,  


-13'd173,  -13'd636,  -13'd598,  13'd293,  13'd73,  -13'd1254,  
13'd271,  -13'd177,  13'd97,  13'd314,  -13'd256,  -13'd914,  
13'd87,  13'd491,  -13'd47,  13'd888,  13'd707,  -13'd979,  
-13'd217,  13'd22,  -13'd683,  13'd80,  -13'd641,  -13'd674,  
13'd267,  -13'd214,  -13'd111,  13'd679,  13'd451,  13'd828,  
13'd911,  13'd295,  -13'd450,  -13'd82,  13'd740,  -13'd327,  
-13'd591,  13'd647,  13'd422,  13'd191,  13'd74,  -13'd474,  
-13'd702,  -13'd46,  13'd374,  13'd417,  -13'd15,  13'd217,  
13'd401,  13'd985,  -13'd866,  -13'd293,  -13'd97,  -13'd80,  
-13'd334,  13'd157,  -13'd24,  -13'd595,  13'd764,  -13'd212,  
13'd305,  -13'd292,  13'd7,  13'd698,  -13'd845,  -13'd367,  
13'd529,  -13'd64,  13'd47,  13'd431,  13'd928,  13'd279,  
13'd3,  13'd837,  13'd733,  13'd536,  13'd313,  13'd264,  
13'd112,  13'd450,  13'd103,  13'd781,  -13'd94,  13'd693,  
-13'd525,  -13'd826,  13'd146,  13'd305,  -13'd1412,  13'd563,  
13'd60,  -13'd27,  13'd292,  13'd347,  13'd131,  13'd604,  

-13'd63,  13'd560,  13'd148,  13'd99,  13'd512,  -13'd813,  
-13'd646,  13'd150,  13'd846,  -13'd438,  -13'd45,  13'd1201,  
-13'd1096,  -13'd95,  -13'd130,  -13'd420,  -13'd345,  -13'd125,  
13'd482,  13'd133,  -13'd100,  13'd1111,  -13'd64,  -13'd541,  
13'd806,  13'd85,  13'd165,  -13'd434,  13'd247,  13'd352,  
-13'd898,  -13'd158,  -13'd504,  13'd711,  13'd207,  13'd351,  
13'd196,  13'd713,  13'd637,  -13'd66,  -13'd1271,  13'd658,  
13'd114,  -13'd71,  -13'd769,  13'd923,  -13'd324,  -13'd407,  
-13'd507,  -13'd16,  13'd684,  -13'd831,  -13'd304,  -13'd33,  
-13'd63,  13'd387,  13'd592,  -13'd161,  13'd1030,  -13'd414,  
-13'd23,  -13'd26,  -13'd325,  13'd361,  -13'd332,  -13'd25,  
13'd270,  13'd441,  -13'd487,  13'd146,  13'd621,  13'd194,  
-13'd282,  -13'd349,  13'd412,  13'd859,  13'd142,  13'd385,  
13'd207,  13'd263,  13'd287,  -13'd650,  13'd521,  13'd441,  
-13'd518,  13'd337,  -13'd676,  13'd222,  -13'd697,  -13'd422,  
13'd434,  -13'd254,  13'd183,  -13'd534,  13'd172,  13'd607,  

-13'd325,  13'd322,  13'd179,  13'd113,  13'd429,  -13'd67,  
-13'd624,  -13'd338,  -13'd11,  -13'd357,  -13'd27,  13'd1115,  
-13'd505,  13'd226,  -13'd276,  13'd218,  -13'd553,  -13'd395,  
13'd596,  13'd34,  13'd416,  13'd482,  13'd258,  -13'd1176,  
13'd620,  -13'd579,  -13'd305,  13'd250,  13'd135,  13'd200,  
-13'd785,  13'd124,  13'd271,  13'd552,  -13'd398,  -13'd686,  
13'd460,  -13'd442,  13'd1082,  13'd128,  -13'd741,  13'd466,  
13'd426,  13'd13,  -13'd533,  13'd632,  -13'd693,  -13'd280,  
-13'd131,  -13'd638,  -13'd401,  -13'd347,  -13'd632,  13'd275,  
13'd15,  -13'd11,  13'd259,  -13'd14,  13'd537,  -13'd117,  
13'd312,  13'd430,  -13'd482,  13'd523,  13'd396,  13'd346,  
13'd438,  13'd237,  -13'd266,  -13'd18,  -13'd497,  13'd390,  
13'd632,  13'd415,  -13'd241,  13'd687,  13'd116,  13'd67,  
-13'd681,  13'd97,  -13'd567,  -13'd106,  -13'd998,  -13'd653,  
13'd526,  13'd1184,  13'd174,  13'd298,  -13'd1242,  13'd299,  
13'd315,  -13'd811,  13'd280,  13'd95,  13'd17,  13'd580,  

-13'd1148,  13'd1061,  13'd1033,  13'd497,  -13'd667,  13'd1113,  
13'd104,  -13'd450,  -13'd457,  -13'd132,  -13'd1040,  13'd297,  
13'd69,  13'd565,  13'd523,  13'd1108,  -13'd1317,  13'd290,  
13'd603,  13'd417,  13'd139,  13'd809,  13'd946,  -13'd615,  
-13'd527,  13'd93,  -13'd477,  -13'd790,  13'd708,  13'd812,  
13'd758,  13'd759,  13'd306,  13'd448,  -13'd389,  -13'd1028,  
13'd138,  -13'd1107,  -13'd184,  -13'd121,  -13'd489,  13'd373,  
13'd154,  13'd407,  13'd299,  13'd754,  13'd726,  13'd130,  
13'd453,  -13'd129,  -13'd462,  -13'd67,  13'd804,  13'd55,  
13'd687,  -13'd472,  -13'd631,  13'd698,  13'd60,  -13'd1275,  
13'd493,  -13'd717,  13'd414,  13'd195,  13'd432,  13'd797,  
13'd258,  13'd83,  13'd571,  -13'd326,  -13'd490,  13'd410,  
13'd885,  13'd185,  13'd260,  13'd819,  13'd115,  -13'd353,  
-13'd901,  13'd160,  -13'd222,  13'd548,  -13'd1192,  13'd944,  
13'd873,  13'd40,  13'd757,  -13'd99,  -13'd15,  -13'd842,  
13'd569,  -13'd335,  13'd300,  -13'd377,  -13'd566,  -13'd1056,  

13'd766,  -13'd267,  13'd392,  13'd145,  -13'd1587,  13'd1301,  
13'd2,  -13'd65,  -13'd528,  13'd206,  -13'd398,  13'd450,  
13'd440,  13'd73,  -13'd440,  -13'd71,  -13'd1061,  13'd30,  
13'd625,  13'd866,  13'd543,  13'd139,  13'd796,  13'd190,  
-13'd265,  -13'd194,  -13'd48,  -13'd539,  13'd271,  13'd623,  
13'd434,  13'd385,  -13'd214,  13'd894,  -13'd599,  13'd60,  
13'd241,  13'd304,  -13'd1184,  -13'd706,  -13'd1129,  -13'd944,  
13'd210,  13'd658,  -13'd531,  13'd900,  13'd371,  13'd173,  
13'd588,  13'd581,  -13'd498,  13'd377,  13'd571,  13'd192,  
13'd1027,  -13'd318,  -13'd43,  13'd261,  13'd543,  -13'd560,  
13'd42,  -13'd563,  13'd272,  -13'd529,  -13'd1468,  13'd608,  
-13'd484,  13'd475,  13'd1371,  -13'd769,  -13'd401,  13'd1757,  
13'd102,  13'd363,  13'd585,  13'd151,  13'd415,  13'd271,  
-13'd94,  13'd554,  13'd292,  13'd853,  -13'd1170,  13'd467,  
-13'd53,  13'd172,  13'd14,  13'd11,  13'd91,  -13'd658,  
13'd873,  -13'd106,  13'd171,  -13'd318,  -13'd669,  13'd349,  


13'd500,  13'd471,  13'd66,  -13'd144,  13'd864,  -13'd465,  
-13'd94,  13'd355,  13'd476,  -13'd384,  -13'd45,  13'd590,  
13'd610,  13'd734,  13'd422,  13'd354,  13'd622,  -13'd838,  
13'd107,  13'd285,  13'd486,  13'd795,  13'd342,  -13'd511,  
-13'd800,  -13'd631,  13'd176,  -13'd200,  -13'd964,  13'd93,  
13'd315,  13'd509,  -13'd342,  13'd718,  -13'd30,  13'd125,  
-13'd1155,  13'd585,  13'd988,  13'd639,  -13'd744,  13'd158,  
-13'd114,  -13'd603,  13'd398,  13'd319,  -13'd683,  13'd289,  
13'd217,  13'd807,  13'd826,  13'd85,  -13'd460,  13'd1309,  
13'd665,  13'd562,  -13'd681,  -13'd88,  13'd517,  13'd249,  
-13'd986,  -13'd28,  -13'd667,  13'd693,  -13'd711,  13'd434,  
-13'd72,  -13'd420,  -13'd514,  13'd12,  13'd403,  13'd344,  
-13'd184,  -13'd374,  13'd47,  13'd662,  13'd263,  13'd478,  
-13'd121,  13'd66,  -13'd269,  -13'd167,  -13'd112,  13'd99,  
13'd429,  -13'd642,  13'd199,  -13'd422,  -13'd896,  -13'd59,  
13'd74,  -13'd416,  -13'd531,  -13'd333,  -13'd357,  -13'd31,  

-13'd796,  13'd812,  13'd786,  13'd109,  13'd406,  13'd836,  
-13'd580,  13'd535,  13'd1333,  -13'd226,  -13'd505,  13'd671,  
13'd208,  -13'd92,  -13'd202,  -13'd55,  13'd299,  -13'd972,  
13'd200,  -13'd57,  -13'd417,  13'd266,  13'd217,  -13'd463,  
-13'd244,  -13'd81,  13'd53,  13'd25,  13'd41,  13'd58,  
-13'd966,  13'd253,  13'd326,  13'd207,  -13'd339,  13'd30,  
-13'd35,  -13'd216,  13'd393,  13'd365,  -13'd1002,  -13'd72,  
-13'd811,  -13'd523,  -13'd139,  -13'd31,  -13'd1777,  13'd44,  
-13'd615,  13'd482,  13'd542,  -13'd460,  -13'd268,  13'd617,  
13'd18,  13'd439,  13'd359,  13'd554,  13'd631,  13'd319,  
-13'd565,  13'd121,  -13'd126,  -13'd316,  13'd139,  13'd148,  
-13'd149,  13'd263,  13'd118,  -13'd30,  13'd346,  13'd7,  
13'd969,  -13'd679,  -13'd280,  -13'd280,  -13'd163,  13'd70,  
13'd219,  13'd287,  13'd383,  -13'd416,  13'd224,  13'd768,  
13'd725,  13'd549,  -13'd596,  -13'd37,  -13'd651,  -13'd77,  
13'd197,  -13'd139,  13'd225,  -13'd384,  13'd201,  -13'd305,  

-13'd862,  -13'd38,  -13'd159,  13'd469,  -13'd624,  13'd438,  
13'd271,  -13'd522,  13'd340,  -13'd862,  -13'd1408,  13'd464,  
-13'd727,  13'd249,  -13'd317,  13'd123,  -13'd651,  -13'd523,  
13'd508,  13'd234,  -13'd119,  13'd327,  -13'd168,  -13'd659,  
13'd564,  13'd152,  13'd781,  -13'd1,  13'd22,  -13'd50,  
-13'd914,  -13'd222,  -13'd413,  -13'd849,  -13'd362,  13'd866,  
13'd899,  -13'd418,  -13'd166,  13'd152,  -13'd1171,  13'd97,  
-13'd431,  -13'd729,  -13'd361,  13'd487,  -13'd519,  -13'd746,  
13'd123,  -13'd1219,  -13'd461,  -13'd523,  -13'd826,  13'd504,  
13'd484,  -13'd426,  -13'd200,  -13'd324,  -13'd133,  -13'd658,  
-13'd499,  -13'd198,  -13'd48,  13'd551,  13'd506,  -13'd766,  
13'd195,  13'd294,  13'd488,  -13'd528,  13'd413,  13'd268,  
13'd432,  -13'd69,  -13'd962,  13'd721,  13'd42,  -13'd213,  
-13'd290,  -13'd468,  -13'd220,  -13'd683,  -13'd254,  -13'd177,  
13'd139,  13'd651,  13'd6,  13'd1148,  -13'd591,  -13'd489,  
-13'd246,  13'd21,  -13'd556,  -13'd756,  13'd363,  -13'd910,  

13'd60,  -13'd216,  -13'd688,  13'd112,  -13'd2177,  -13'd519,  
-13'd343,  -13'd363,  -13'd765,  -13'd171,  -13'd1544,  -13'd346,  
-13'd534,  13'd4,  13'd404,  13'd411,  -13'd1656,  13'd536,  
-13'd70,  -13'd372,  -13'd535,  13'd717,  13'd588,  -13'd273,  
13'd359,  13'd744,  -13'd244,  13'd71,  13'd859,  -13'd989,  
13'd462,  -13'd564,  -13'd378,  13'd367,  -13'd1320,  -13'd321,  
13'd137,  -13'd426,  -13'd1076,  -13'd746,  -13'd342,  -13'd891,  
13'd771,  -13'd122,  -13'd525,  13'd156,  -13'd306,  -13'd1207,  
13'd1129,  13'd620,  -13'd462,  -13'd570,  -13'd203,  -13'd501,  
-13'd75,  13'd102,  -13'd180,  -13'd76,  13'd243,  -13'd978,  
-13'd374,  -13'd1312,  -13'd930,  -13'd479,  -13'd48,  -13'd452,  
-13'd522,  -13'd196,  13'd458,  13'd641,  -13'd426,  13'd515,  
-13'd221,  -13'd439,  -13'd476,  13'd872,  13'd488,  -13'd1117,  
-13'd488,  13'd40,  13'd191,  13'd33,  -13'd1139,  13'd643,  
13'd432,  13'd225,  -13'd231,  13'd743,  13'd325,  -13'd189,  
-13'd661,  13'd227,  -13'd74,  -13'd179,  -13'd319,  13'd202,  

-13'd181,  13'd91,  -13'd114,  13'd278,  -13'd738,  13'd256,  
13'd258,  13'd742,  13'd189,  13'd79,  -13'd751,  13'd976,  
13'd530,  -13'd97,  13'd259,  13'd249,  -13'd457,  -13'd600,  
13'd1090,  13'd251,  13'd48,  13'd198,  13'd512,  -13'd260,  
13'd270,  13'd160,  13'd145,  -13'd126,  13'd238,  -13'd283,  
13'd597,  -13'd50,  13'd241,  13'd997,  -13'd60,  -13'd973,  
-13'd44,  13'd543,  -13'd249,  -13'd678,  -13'd87,  -13'd49,  
13'd771,  13'd197,  -13'd147,  13'd510,  13'd770,  -13'd1073,  
13'd1242,  -13'd402,  -13'd932,  -13'd154,  13'd1106,  -13'd32,  
13'd168,  -13'd27,  -13'd550,  13'd327,  -13'd790,  -13'd729,  
-13'd558,  -13'd459,  -13'd1301,  -13'd1100,  13'd255,  -13'd623,  
-13'd608,  13'd68,  -13'd82,  13'd287,  -13'd1665,  13'd1256,  
13'd113,  -13'd95,  -13'd65,  -13'd501,  13'd667,  -13'd337,  
13'd658,  -13'd313,  13'd768,  13'd653,  -13'd935,  13'd138,  
13'd749,  13'd34,  13'd77,  13'd684,  -13'd33,  -13'd61,  
13'd12,  -13'd355,  13'd187,  13'd361,  -13'd718,  13'd908,  


-13'd251,  13'd25,  -13'd335,  -13'd951,  13'd556,  13'd946,  
-13'd912,  13'd360,  -13'd104,  -13'd88,  -13'd273,  -13'd65,  
13'd1076,  -13'd356,  -13'd378,  13'd203,  -13'd133,  -13'd305,  
-13'd710,  -13'd635,  13'd208,  -13'd79,  -13'd377,  -13'd276,  
13'd337,  13'd282,  -13'd211,  -13'd720,  13'd81,  -13'd323,  
-13'd749,  13'd781,  13'd441,  -13'd173,  -13'd554,  13'd461,  
-13'd114,  13'd677,  13'd1104,  13'd162,  -13'd609,  13'd34,  
-13'd470,  -13'd775,  13'd455,  13'd135,  13'd440,  -13'd987,  
-13'd706,  13'd1328,  13'd1515,  13'd857,  -13'd1538,  13'd894,  
13'd771,  -13'd455,  13'd279,  13'd202,  -13'd304,  13'd49,  
-13'd580,  13'd387,  13'd164,  -13'd131,  -13'd313,  13'd566,  
-13'd661,  13'd287,  -13'd718,  -13'd154,  -13'd683,  13'd213,  
13'd226,  -13'd503,  -13'd1101,  -13'd824,  13'd352,  -13'd279,  
-13'd137,  13'd638,  13'd572,  13'd264,  -13'd585,  -13'd73,  
-13'd123,  -13'd228,  -13'd340,  -13'd110,  -13'd820,  -13'd153,  
13'd156,  -13'd249,  -13'd651,  -13'd612,  13'd705,  -13'd10,  

-13'd560,  13'd196,  13'd565,  -13'd250,  -13'd832,  13'd338,  
-13'd706,  13'd504,  13'd386,  -13'd174,  -13'd1434,  13'd784,  
13'd219,  13'd359,  13'd404,  -13'd56,  13'd184,  -13'd811,  
-13'd315,  -13'd1068,  -13'd230,  13'd178,  -13'd984,  13'd485,  
-13'd154,  -13'd118,  -13'd65,  -13'd531,  13'd24,  13'd953,  
-13'd174,  13'd115,  13'd34,  -13'd129,  -13'd332,  13'd543,  
13'd558,  13'd318,  -13'd46,  13'd183,  -13'd1154,  13'd819,  
-13'd964,  -13'd147,  -13'd815,  -13'd422,  -13'd454,  -13'd16,  
13'd601,  13'd625,  13'd925,  13'd577,  -13'd1465,  13'd1087,  
13'd859,  13'd118,  -13'd543,  13'd532,  13'd486,  -13'd1167,  
13'd193,  -13'd1000,  -13'd785,  -13'd543,  13'd1019,  -13'd86,  
-13'd34,  13'd404,  13'd87,  -13'd243,  -13'd287,  -13'd26,  
-13'd27,  -13'd765,  -13'd386,  -13'd309,  13'd1112,  -13'd347,  
-13'd350,  -13'd138,  13'd858,  13'd98,  -13'd314,  -13'd59,  
-13'd630,  13'd135,  -13'd231,  -13'd1037,  -13'd463,  -13'd403,  
13'd485,  13'd169,  -13'd218,  -13'd71,  13'd781,  -13'd415,  

-13'd547,  13'd473,  -13'd247,  13'd526,  -13'd1578,  13'd93,  
13'd865,  -13'd838,  -13'd393,  13'd152,  -13'd398,  13'd152,  
-13'd251,  13'd660,  -13'd466,  13'd44,  -13'd489,  13'd247,  
-13'd462,  -13'd956,  -13'd532,  13'd384,  -13'd405,  -13'd495,  
-13'd622,  13'd386,  13'd313,  -13'd42,  -13'd212,  13'd134,  
-13'd420,  -13'd1213,  13'd167,  -13'd235,  -13'd590,  13'd150,  
13'd314,  -13'd744,  -13'd286,  -13'd60,  -13'd560,  -13'd534,  
-13'd438,  -13'd458,  13'd351,  -13'd237,  -13'd15,  -13'd226,  
13'd683,  13'd349,  -13'd381,  13'd221,  -13'd161,  -13'd268,  
13'd448,  13'd679,  -13'd607,  -13'd274,  13'd201,  -13'd1081,  
-13'd711,  13'd144,  -13'd1130,  -13'd597,  13'd221,  -13'd1589,  
-13'd785,  13'd14,  13'd307,  13'd508,  -13'd473,  13'd970,  
-13'd390,  13'd88,  -13'd487,  -13'd350,  13'd600,  -13'd66,  
-13'd244,  13'd125,  13'd401,  -13'd342,  13'd609,  -13'd375,  
-13'd212,  -13'd567,  -13'd280,  13'd66,  -13'd774,  -13'd868,  
-13'd131,  13'd271,  -13'd230,  -13'd648,  13'd500,  13'd976,  

13'd718,  -13'd480,  -13'd608,  13'd330,  -13'd875,  -13'd426,  
-13'd89,  13'd45,  13'd416,  -13'd315,  -13'd311,  13'd370,  
13'd155,  13'd197,  13'd290,  13'd200,  -13'd925,  13'd994,  
-13'd782,  -13'd998,  -13'd872,  -13'd202,  -13'd885,  -13'd847,  
13'd263,  13'd15,  13'd595,  -13'd119,  -13'd154,  -13'd229,  
13'd95,  -13'd66,  -13'd354,  -13'd86,  -13'd131,  -13'd842,  
13'd22,  13'd301,  -13'd493,  13'd185,  13'd778,  -13'd752,  
-13'd634,  -13'd582,  13'd95,  -13'd511,  -13'd228,  13'd173,  
-13'd744,  -13'd85,  -13'd609,  -13'd964,  13'd87,  13'd235,  
13'd367,  13'd587,  -13'd311,  13'd60,  13'd1274,  13'd202,  
-13'd525,  -13'd626,  -13'd806,  -13'd1234,  13'd366,  -13'd882,  
13'd172,  -13'd1002,  -13'd250,  13'd211,  13'd68,  13'd233,  
-13'd1224,  -13'd360,  -13'd16,  -13'd929,  -13'd94,  -13'd408,  
13'd238,  13'd618,  13'd737,  -13'd12,  -13'd618,  13'd81,  
13'd544,  13'd38,  -13'd481,  13'd238,  -13'd413,  -13'd106,  
-13'd866,  13'd183,  13'd502,  -13'd192,  -13'd309,  13'd9,  

-13'd144,  -13'd489,  -13'd978,  13'd462,  -13'd447,  -13'd721,  
-13'd411,  -13'd28,  13'd911,  13'd413,  -13'd580,  13'd946,  
13'd692,  -13'd725,  -13'd533,  13'd744,  -13'd272,  13'd63,  
-13'd200,  -13'd465,  -13'd196,  -13'd412,  -13'd465,  -13'd878,  
13'd225,  -13'd127,  -13'd177,  13'd77,  -13'd83,  -13'd58,  
-13'd83,  -13'd813,  -13'd487,  -13'd282,  -13'd913,  -13'd188,  
13'd374,  13'd988,  -13'd150,  -13'd100,  13'd316,  13'd287,  
-13'd703,  -13'd433,  -13'd506,  -13'd276,  -13'd62,  13'd346,  
13'd488,  -13'd955,  -13'd294,  -13'd265,  13'd18,  -13'd98,  
-13'd5,  -13'd496,  13'd301,  -13'd499,  13'd203,  -13'd805,  
-13'd806,  13'd857,  -13'd216,  -13'd672,  13'd274,  -13'd555,  
-13'd95,  -13'd46,  -13'd81,  13'd137,  13'd210,  -13'd1397,  
-13'd1323,  -13'd600,  13'd131,  -13'd936,  -13'd988,  13'd542,  
13'd871,  13'd645,  -13'd170,  13'd104,  -13'd698,  -13'd158,  
13'd436,  -13'd1003,  13'd217,  -13'd33,  -13'd339,  -13'd289,  
-13'd183,  -13'd218,  -13'd42,  13'd426,  -13'd637,  13'd99
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule


module bias_fc1_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC1-1][0:`OUTPUT_NUM_FC1-1][`WD_BIAS:0] weight	 = {
-24'd219560,  -24'd253697,  -24'd55433,  -24'd97677,  24'd293697,  -24'd243881,  24'd320084,  24'd224550,  24'd239030,  24'd511222,  24'd91710,  24'd236129,  24'd189478,  24'd189715,  24'd237750,  24'd85050,  
24'd84279,  -24'd41102,  24'd389770,  24'd141391,  -24'd114359,  24'd179309,  24'd335280,  24'd91496,  -24'd304524,  24'd51767,  24'd50531,  24'd398249,  24'd125193,  24'd59246,  24'd302096,  -24'd391546,  
-24'd8719,  -24'd143200,  24'd86710,  -24'd121286,  -24'd17574,  24'd193986,  24'd334251,  24'd418338,  -24'd29725,  -24'd164781,  24'd19566,  24'd369659,  24'd369117,  24'd485986,  24'd255667,  24'd184972,  
-24'd350874,  24'd83616,  -24'd113753,  24'd50318,  -24'd218172,  24'd245365,  -24'd212866,  -24'd167942,  24'd24266,  -24'd290894,  -24'd45370,  24'd333035,  24'd76391,  24'd331919,  24'd249570,  24'd116175,  
24'd314113,  24'd322302,  -24'd387295,  -24'd139803,  24'd555959,  24'd41557,  -24'd71756,  24'd250106,  24'd125286,  24'd209370,  -24'd167080,  24'd330490,  24'd186924,  24'd87729,  -24'd220844,  24'd340936,  
-24'd135930,  24'd117423,  24'd224274,  -24'd3834,  -24'd49645,  -24'd105418,  24'd52762,  24'd96732,  -24'd152523,  24'd141711,  24'd257837,  -24'd91013,  24'd178395,  24'd55568,  -24'd93767,  -24'd131308,  
24'd155983,  -24'd449369,  24'd184192,  -24'd39257,  -24'd140313,  24'd360847,  24'd255272,  24'd73788,  -24'd213748,  24'd163158,  24'd149546,  24'd206663,  -24'd58642,  -24'd77157,  -24'd41775,  24'd140758,  
24'd396969,  24'd190957,  24'd87027,  -24'd48891,  24'd157309,  -24'd282668,  -24'd283377,  -24'd195665
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_fc1_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1*`OUTPUT_BATCH_FC1)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV2*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC1*`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1-1][0:`OUTPUT_NUM_FC1-1][0:`OUTPUT_NUM_CONV2-1][`WD:0] weight	 = {
-13'd176,  13'd98,  -13'd104,  13'd1000,  -13'd8,  13'd1,  13'd241,  -13'd876,  13'd448,  13'd278,  -13'd141,  -13'd266,  13'd411,  -13'd460,  -13'd356,  -13'd96,  
13'd879,  13'd93,  13'd480,  13'd423,  -13'd435,  13'd331,  -13'd577,  13'd490,  13'd85,  -13'd59,  13'd8,  13'd131,  13'd504,  -13'd281,  -13'd27,  13'd152,  
13'd322,  -13'd557,  13'd170,  -13'd505,  -13'd676,  -13'd311,  13'd85,  -13'd574,  13'd242,  -13'd470,  13'd858,  13'd512,  13'd630,  -13'd293,  -13'd440,  13'd990,  
13'd240,  13'd106,  13'd366,  13'd1,  -13'd401,  13'd669,  13'd858,  13'd286,  13'd642,  -13'd16,  13'd570,  13'd7,  13'd351,  13'd705,  -13'd222,  -13'd87,  
13'd917,  13'd819,  -13'd656,  13'd320,  13'd938,  13'd673,  13'd648,  13'd579,  13'd391,  -13'd260,  13'd92,  13'd659,  13'd914,  13'd350,  -13'd1016,  13'd264,  
13'd515,  13'd340,  -13'd509,  13'd372,  13'd422,  -13'd170,  13'd386,  -13'd807,  -13'd279,  -13'd401,  13'd1053,  -13'd232,  -13'd68,  -13'd459,  13'd764,  -13'd26,  
13'd81,  13'd267,  -13'd297,  -13'd337,  -13'd72,  13'd393,  13'd195,  -13'd28,  13'd292,  13'd182,  13'd865,  13'd243,  -13'd576,  -13'd302,  -13'd951,  -13'd710,  
13'd167,  -13'd532,  -13'd280,  -13'd447,  -13'd50,  13'd213,  13'd102,  -13'd496,  13'd136,  13'd698,  -13'd100,  13'd238,  13'd835,  -13'd97,  -13'd368,  13'd298,  
13'd563,  -13'd671,  -13'd480,  -13'd666,  -13'd43,  13'd126,  -13'd315,  -13'd617,  -13'd574,  -13'd883,  -13'd376,  -13'd341,  13'd530,  13'd716,  13'd297,  13'd223,  
-13'd179,  -13'd72,  -13'd1505,  -13'd297,  -13'd417,  -13'd223,  -13'd46,  -13'd100,  -13'd534,  -13'd602,  13'd349,  -13'd427,  -13'd365,  -13'd373,  13'd372,  -13'd645,  
-13'd185,  13'd70,  13'd823,  -13'd880,  -13'd223,  -13'd507,  -13'd98,  -13'd479,  -13'd243,  -13'd521,  -13'd614,  13'd276,  13'd323,  -13'd112,  -13'd26,  -13'd80,  
-13'd50,  13'd675,  13'd443,  -13'd706,  -13'd566,  13'd12,  13'd434,  -13'd193,  13'd294,  13'd253,  -13'd656,  -13'd124,  -13'd609,  13'd720,  -13'd522,  -13'd218,  
-13'd4,  -13'd329,  -13'd448,  -13'd608,  -13'd411,  -13'd534,  -13'd570,  -13'd717,  -13'd606,  -13'd351,  -13'd950,  -13'd410,  13'd176,  13'd765,  -13'd343,  -13'd266,  
13'd8,  -13'd327,  13'd614,  13'd392,  -13'd7,  -13'd1316,  -13'd231,  -13'd228,  13'd39,  13'd461,  -13'd740,  -13'd469,  13'd36,  13'd473,  -13'd542,  -13'd12,  
-13'd1086,  -13'd686,  13'd281,  13'd351,  -13'd120,  -13'd934,  13'd77,  -13'd760,  -13'd7,  13'd790,  -13'd57,  13'd403,  -13'd509,  -13'd225,  -13'd11,  -13'd998,  
-13'd251,  -13'd332,  13'd135,  13'd672,  13'd477,  -13'd69,  -13'd1154,  -13'd149,  13'd336,  -13'd14,  -13'd641,  -13'd629,  13'd205,  -13'd31,  13'd904,  -13'd123,  
-13'd432,  -13'd732,  -13'd144,  13'd1202,  13'd394,  -13'd103,  -13'd324,  13'd372,  -13'd387,  -13'd29,  13'd832,  -13'd552,  -13'd78,  -13'd234,  -13'd133,  -13'd690,  
13'd37,  -13'd104,  13'd223,  13'd92,  -13'd187,  -13'd801,  -13'd1365,  13'd76,  -13'd1211,  13'd684,  -13'd110,  -13'd395,  13'd393,  13'd5,  -13'd171,  13'd681,  
-13'd123,  -13'd486,  13'd233,  13'd367,  -13'd709,  13'd77,  13'd98,  -13'd30,  -13'd336,  -13'd668,  -13'd622,  13'd687,  13'd656,  -13'd10,  13'd135,  13'd450,  
-13'd341,  -13'd471,  -13'd377,  -13'd283,  -13'd193,  -13'd112,  13'd582,  13'd152,  13'd557,  -13'd485,  13'd71,  13'd811,  -13'd161,  -13'd149,  -13'd17,  -13'd275,  
-13'd522,  13'd735,  -13'd552,  -13'd412,  13'd108,  13'd288,  -13'd535,  13'd362,  13'd1378,  13'd187,  13'd1088,  -13'd798,  -13'd25,  -13'd667,  13'd66,  -13'd15,  
-13'd421,  13'd154,  -13'd1037,  -13'd384,  -13'd297,  -13'd417,  -13'd1162,  -13'd667,  13'd627,  -13'd743,  13'd393,  13'd44,  -13'd112,  -13'd1157,  13'd53,  13'd580,  
13'd69,  -13'd101,  -13'd732,  13'd91,  -13'd1161,  -13'd556,  -13'd872,  13'd351,  -13'd338,  -13'd241,  13'd430,  -13'd122,  -13'd234,  13'd800,  13'd153,  -13'd60,  
-13'd436,  13'd71,  13'd983,  -13'd650,  -13'd736,  -13'd16,  13'd745,  -13'd440,  13'd18,  -13'd181,  -13'd380,  13'd169,  13'd160,  13'd1173,  13'd823,  13'd411,  
13'd665,  13'd228,  13'd657,  13'd476,  -13'd5,  13'd327,  13'd672,  13'd130,  13'd120,  -13'd1123,  -13'd349,  13'd420,  -13'd249,  -13'd236,  13'd460,  13'd492,  

-13'd212,  -13'd3,  -13'd132,  13'd240,  -13'd277,  13'd402,  -13'd555,  -13'd103,  -13'd762,  -13'd175,  13'd51,  13'd289,  -13'd87,  -13'd207,  13'd206,  13'd374,  
-13'd625,  -13'd682,  -13'd377,  -13'd412,  -13'd612,  -13'd465,  -13'd54,  -13'd108,  13'd56,  -13'd504,  13'd165,  13'd533,  13'd554,  13'd203,  -13'd873,  -13'd422,  
-13'd228,  -13'd418,  -13'd246,  -13'd346,  -13'd113,  13'd541,  -13'd236,  13'd343,  13'd217,  -13'd637,  -13'd210,  -13'd385,  -13'd111,  13'd182,  13'd244,  -13'd460,  
13'd274,  13'd375,  -13'd73,  13'd195,  -13'd256,  -13'd58,  -13'd851,  -13'd317,  -13'd462,  -13'd156,  -13'd890,  -13'd113,  -13'd328,  -13'd254,  13'd10,  13'd15,  
13'd702,  -13'd277,  -13'd170,  -13'd454,  13'd264,  -13'd852,  -13'd305,  -13'd172,  -13'd357,  13'd222,  -13'd829,  -13'd39,  13'd168,  13'd139,  -13'd66,  -13'd779,  
13'd127,  13'd23,  13'd548,  -13'd411,  13'd176,  13'd372,  -13'd314,  -13'd479,  -13'd227,  13'd479,  -13'd549,  13'd202,  13'd706,  13'd69,  -13'd265,  -13'd774,  
-13'd111,  -13'd200,  -13'd500,  -13'd157,  -13'd126,  -13'd178,  13'd237,  -13'd352,  -13'd527,  13'd534,  13'd320,  -13'd657,  -13'd21,  13'd244,  -13'd135,  -13'd537,  
13'd472,  -13'd425,  13'd169,  13'd375,  13'd411,  13'd381,  -13'd544,  13'd158,  13'd214,  13'd144,  -13'd141,  13'd311,  -13'd189,  -13'd143,  13'd373,  13'd341,  
-13'd21,  -13'd605,  13'd18,  -13'd469,  -13'd176,  13'd160,  13'd382,  -13'd460,  13'd99,  -13'd81,  -13'd70,  -13'd532,  -13'd993,  -13'd390,  13'd22,  -13'd918,  
13'd104,  -13'd134,  -13'd144,  -13'd397,  13'd185,  13'd63,  -13'd450,  -13'd139,  13'd157,  13'd121,  -13'd19,  -13'd99,  13'd46,  -13'd170,  -13'd778,  -13'd590,  
-13'd259,  -13'd254,  -13'd32,  -13'd788,  -13'd729,  -13'd182,  -13'd533,  -13'd9,  -13'd802,  13'd128,  13'd143,  -13'd303,  -13'd418,  13'd18,  -13'd156,  -13'd37,  
-13'd814,  -13'd758,  -13'd36,  -13'd280,  13'd312,  -13'd550,  13'd71,  -13'd125,  13'd214,  13'd577,  13'd103,  -13'd398,  13'd217,  -13'd146,  -13'd34,  13'd77,  
13'd104,  13'd44,  -13'd724,  13'd374,  13'd340,  -13'd545,  13'd63,  -13'd398,  13'd284,  -13'd339,  13'd257,  13'd551,  13'd228,  -13'd443,  13'd252,  -13'd466,  
-13'd86,  -13'd145,  -13'd373,  13'd548,  -13'd639,  13'd459,  13'd198,  -13'd228,  -13'd254,  -13'd819,  -13'd471,  -13'd412,  13'd168,  13'd259,  -13'd387,  13'd137,  
-13'd196,  -13'd134,  13'd93,  -13'd408,  13'd380,  -13'd149,  -13'd681,  13'd298,  -13'd188,  -13'd117,  -13'd279,  -13'd293,  -13'd249,  -13'd318,  -13'd470,  -13'd259,  
13'd591,  13'd188,  -13'd422,  -13'd420,  -13'd392,  -13'd240,  -13'd757,  -13'd471,  13'd402,  -13'd427,  -13'd671,  13'd44,  -13'd50,  -13'd304,  -13'd342,  -13'd383,  
-13'd808,  13'd269,  -13'd59,  13'd260,  -13'd377,  13'd190,  13'd175,  -13'd113,  -13'd739,  13'd172,  -13'd294,  -13'd601,  -13'd788,  -13'd325,  -13'd532,  13'd522,  
13'd134,  13'd482,  13'd21,  13'd377,  13'd515,  -13'd300,  13'd322,  -13'd310,  -13'd519,  13'd41,  -13'd376,  13'd495,  -13'd10,  -13'd241,  13'd227,  -13'd538,  
-13'd78,  -13'd224,  -13'd127,  -13'd321,  -13'd385,  13'd88,  -13'd509,  -13'd203,  13'd69,  13'd226,  -13'd370,  -13'd535,  -13'd700,  -13'd189,  -13'd274,  -13'd362,  
13'd110,  -13'd459,  -13'd29,  -13'd268,  -13'd494,  -13'd435,  -13'd2,  -13'd766,  -13'd50,  -13'd226,  -13'd562,  13'd363,  13'd143,  -13'd586,  13'd196,  13'd20,  
-13'd419,  13'd146,  13'd288,  -13'd491,  -13'd697,  -13'd92,  -13'd639,  13'd93,  -13'd30,  -13'd837,  13'd127,  -13'd185,  -13'd265,  -13'd848,  13'd235,  13'd48,  
13'd374,  -13'd709,  -13'd202,  -13'd154,  -13'd327,  -13'd384,  -13'd158,  13'd43,  13'd597,  -13'd159,  -13'd794,  13'd7,  13'd391,  -13'd581,  -13'd33,  -13'd477,  
13'd91,  -13'd68,  13'd663,  13'd96,  -13'd442,  -13'd194,  13'd456,  13'd124,  13'd139,  13'd482,  13'd93,  -13'd668,  -13'd314,  -13'd52,  -13'd300,  13'd396,  
-13'd359,  -13'd646,  13'd96,  -13'd589,  -13'd102,  13'd458,  -13'd166,  -13'd88,  -13'd248,  -13'd274,  -13'd78,  -13'd82,  -13'd341,  -13'd521,  13'd231,  -13'd85,  
-13'd158,  -13'd492,  13'd92,  13'd643,  -13'd265,  -13'd516,  -13'd694,  -13'd415,  13'd304,  13'd37,  13'd129,  -13'd127,  -13'd43,  -13'd463,  13'd357,  13'd263,  

-13'd435,  -13'd469,  13'd781,  -13'd433,  -13'd501,  13'd261,  -13'd1237,  13'd199,  13'd620,  -13'd549,  -13'd936,  13'd121,  -13'd122,  13'd197,  13'd609,  13'd103,  
13'd125,  -13'd201,  13'd1532,  -13'd186,  -13'd66,  13'd327,  13'd102,  -13'd718,  13'd132,  13'd627,  -13'd1205,  13'd325,  13'd252,  -13'd208,  13'd239,  -13'd364,  
-13'd526,  13'd65,  13'd142,  -13'd601,  13'd533,  13'd170,  13'd710,  -13'd224,  -13'd258,  13'd30,  -13'd31,  13'd507,  -13'd406,  13'd1930,  -13'd139,  -13'd404,  
-13'd473,  13'd482,  13'd472,  13'd444,  -13'd88,  13'd60,  13'd479,  -13'd274,  13'd664,  -13'd22,  -13'd96,  -13'd581,  -13'd626,  13'd952,  13'd267,  -13'd8,  
13'd1006,  13'd1238,  -13'd256,  -13'd224,  -13'd130,  -13'd133,  13'd830,  13'd327,  13'd351,  13'd95,  -13'd349,  13'd109,  -13'd361,  -13'd370,  13'd185,  13'd412,  
13'd3,  13'd96,  13'd836,  13'd650,  13'd519,  13'd213,  -13'd1158,  13'd318,  -13'd672,  13'd464,  -13'd640,  -13'd98,  -13'd232,  13'd527,  -13'd9,  13'd242,  
-13'd185,  13'd494,  13'd28,  -13'd382,  -13'd100,  -13'd98,  13'd333,  13'd351,  13'd26,  13'd212,  13'd83,  -13'd35,  -13'd32,  -13'd408,  13'd269,  -13'd379,  
-13'd438,  -13'd949,  13'd475,  -13'd634,  -13'd804,  -13'd598,  13'd328,  13'd159,  13'd13,  -13'd156,  -13'd813,  -13'd460,  -13'd259,  13'd88,  13'd717,  -13'd68,  
13'd430,  13'd15,  -13'd99,  -13'd185,  -13'd601,  13'd2,  13'd34,  -13'd347,  13'd280,  -13'd543,  -13'd8,  -13'd306,  -13'd52,  13'd694,  -13'd384,  -13'd665,  
13'd1097,  13'd271,  -13'd173,  -13'd273,  -13'd208,  -13'd370,  13'd922,  -13'd241,  13'd637,  -13'd250,  13'd370,  13'd203,  13'd1077,  13'd406,  -13'd263,  13'd364,  
13'd220,  13'd100,  13'd146,  -13'd309,  13'd581,  -13'd257,  -13'd320,  13'd107,  -13'd490,  -13'd600,  13'd0,  13'd245,  -13'd799,  -13'd11,  -13'd73,  13'd156,  
13'd501,  13'd538,  13'd227,  -13'd42,  13'd136,  -13'd47,  -13'd99,  13'd673,  -13'd772,  -13'd250,  13'd51,  -13'd353,  -13'd251,  -13'd20,  13'd57,  -13'd255,  
13'd343,  13'd793,  -13'd589,  -13'd323,  13'd30,  13'd751,  13'd101,  13'd229,  13'd455,  13'd396,  13'd188,  -13'd590,  13'd748,  -13'd753,  -13'd512,  -13'd832,  
13'd101,  -13'd195,  13'd253,  13'd906,  13'd190,  13'd456,  -13'd392,  13'd643,  -13'd204,  -13'd153,  13'd87,  -13'd400,  -13'd42,  13'd206,  13'd187,  -13'd40,  
13'd1315,  13'd791,  -13'd271,  -13'd114,  13'd234,  13'd256,  -13'd437,  -13'd453,  13'd253,  -13'd638,  -13'd290,  13'd93,  13'd964,  -13'd326,  13'd465,  13'd864,  
13'd783,  -13'd564,  -13'd236,  -13'd98,  -13'd525,  -13'd462,  13'd210,  -13'd491,  13'd21,  -13'd492,  -13'd722,  13'd706,  -13'd822,  13'd102,  -13'd354,  13'd30,  
13'd816,  13'd484,  13'd426,  -13'd378,  -13'd282,  13'd109,  13'd333,  -13'd162,  13'd657,  13'd727,  -13'd619,  13'd122,  13'd511,  13'd1129,  -13'd255,  13'd90,  
-13'd271,  -13'd33,  -13'd434,  13'd631,  13'd268,  -13'd141,  13'd216,  13'd45,  13'd525,  -13'd43,  13'd420,  13'd111,  -13'd8,  -13'd203,  -13'd563,  13'd144,  
-13'd797,  13'd128,  -13'd806,  -13'd601,  -13'd12,  -13'd535,  -13'd95,  13'd735,  -13'd874,  13'd747,  -13'd256,  -13'd256,  -13'd1082,  -13'd275,  -13'd345,  13'd362,  
13'd135,  -13'd571,  -13'd487,  -13'd791,  13'd145,  -13'd446,  -13'd280,  -13'd286,  -13'd577,  -13'd348,  -13'd39,  13'd236,  13'd376,  -13'd122,  -13'd759,  13'd59,  
13'd1164,  13'd153,  13'd947,  -13'd410,  -13'd584,  13'd671,  -13'd207,  13'd621,  13'd204,  13'd736,  -13'd4,  13'd647,  13'd81,  13'd1155,  13'd511,  13'd586,  
13'd107,  -13'd239,  13'd711,  13'd304,  13'd84,  -13'd789,  -13'd199,  13'd389,  13'd429,  -13'd332,  13'd162,  13'd610,  13'd201,  13'd354,  -13'd238,  -13'd343,  
-13'd547,  13'd132,  -13'd261,  -13'd183,  -13'd136,  -13'd286,  13'd23,  13'd807,  13'd327,  -13'd314,  13'd277,  13'd178,  -13'd121,  13'd524,  13'd24,  -13'd12,  
-13'd387,  -13'd779,  -13'd385,  -13'd297,  13'd620,  -13'd636,  13'd177,  -13'd422,  -13'd938,  13'd80,  -13'd29,  -13'd36,  -13'd491,  -13'd82,  -13'd905,  -13'd335,  
-13'd836,  -13'd1131,  13'd309,  -13'd158,  -13'd444,  -13'd184,  -13'd286,  -13'd438,  -13'd441,  -13'd742,  -13'd162,  -13'd371,  13'd172,  -13'd175,  -13'd953,  -13'd253,  

-13'd6,  13'd205,  13'd324,  13'd119,  13'd181,  13'd407,  -13'd612,  13'd491,  -13'd243,  13'd552,  -13'd342,  -13'd361,  13'd134,  13'd152,  13'd182,  13'd152,  
13'd367,  -13'd101,  13'd9,  -13'd48,  13'd597,  13'd464,  -13'd606,  13'd15,  -13'd218,  -13'd303,  -13'd594,  -13'd305,  -13'd245,  13'd359,  13'd267,  13'd153,  
13'd283,  -13'd206,  -13'd274,  13'd194,  -13'd137,  -13'd100,  13'd256,  -13'd312,  -13'd158,  -13'd412,  13'd364,  -13'd819,  -13'd628,  -13'd187,  13'd134,  13'd82,  
-13'd556,  -13'd234,  -13'd83,  -13'd678,  -13'd121,  13'd170,  -13'd153,  -13'd147,  -13'd337,  13'd352,  -13'd479,  -13'd434,  -13'd175,  13'd386,  13'd441,  -13'd624,  
13'd341,  -13'd801,  -13'd390,  -13'd451,  -13'd97,  13'd129,  -13'd407,  -13'd382,  13'd113,  13'd214,  13'd261,  -13'd668,  -13'd578,  -13'd54,  -13'd472,  13'd644,  
-13'd432,  -13'd616,  13'd230,  -13'd192,  -13'd353,  13'd19,  -13'd203,  13'd209,  13'd157,  13'd559,  -13'd213,  13'd303,  13'd166,  -13'd539,  -13'd30,  13'd51,  
13'd140,  -13'd18,  -13'd336,  -13'd622,  -13'd741,  13'd682,  13'd35,  13'd48,  -13'd509,  13'd91,  13'd34,  -13'd341,  -13'd157,  -13'd242,  -13'd468,  13'd178,  
-13'd794,  -13'd505,  13'd87,  -13'd597,  -13'd90,  -13'd215,  -13'd456,  13'd287,  13'd26,  -13'd488,  -13'd201,  -13'd215,  -13'd96,  -13'd271,  13'd701,  -13'd207,  
13'd143,  -13'd150,  -13'd224,  -13'd523,  13'd140,  -13'd375,  -13'd633,  -13'd486,  -13'd325,  -13'd573,  13'd718,  -13'd536,  -13'd631,  -13'd256,  -13'd403,  -13'd143,  
-13'd598,  -13'd71,  13'd303,  -13'd355,  -13'd37,  -13'd233,  -13'd687,  13'd621,  -13'd404,  13'd166,  -13'd81,  -13'd538,  -13'd782,  -13'd165,  -13'd651,  13'd15,  
-13'd532,  -13'd31,  13'd63,  -13'd307,  13'd519,  -13'd166,  -13'd307,  -13'd50,  13'd145,  -13'd553,  13'd60,  13'd26,  -13'd597,  13'd669,  -13'd236,  -13'd120,  
-13'd27,  -13'd738,  -13'd329,  -13'd512,  13'd58,  -13'd129,  13'd172,  -13'd583,  13'd455,  -13'd497,  -13'd312,  13'd669,  -13'd314,  -13'd145,  -13'd37,  13'd228,  
-13'd462,  13'd538,  -13'd10,  -13'd335,  13'd262,  13'd188,  13'd160,  13'd151,  -13'd770,  13'd117,  -13'd208,  -13'd262,  13'd136,  -13'd290,  13'd206,  13'd230,  
-13'd102,  13'd72,  -13'd460,  -13'd682,  13'd493,  -13'd154,  -13'd438,  -13'd228,  -13'd16,  -13'd846,  -13'd471,  -13'd365,  -13'd468,  -13'd535,  -13'd330,  13'd441,  
-13'd289,  13'd408,  -13'd433,  13'd647,  13'd424,  -13'd208,  13'd293,  13'd36,  -13'd400,  -13'd280,  13'd457,  13'd97,  -13'd191,  -13'd233,  -13'd309,  13'd211,  
13'd161,  13'd18,  13'd287,  13'd114,  13'd94,  13'd443,  -13'd249,  -13'd207,  -13'd184,  -13'd769,  -13'd206,  -13'd167,  -13'd711,  -13'd464,  13'd177,  13'd613,  
-13'd301,  -13'd90,  -13'd28,  -13'd531,  13'd316,  -13'd192,  -13'd65,  13'd108,  -13'd179,  -13'd183,  13'd449,  -13'd636,  13'd601,  -13'd616,  -13'd458,  13'd703,  
13'd278,  -13'd65,  -13'd433,  13'd116,  -13'd594,  -13'd393,  -13'd351,  13'd191,  13'd76,  -13'd4,  -13'd694,  -13'd393,  -13'd273,  13'd206,  -13'd473,  -13'd217,  
-13'd449,  -13'd2,  -13'd511,  13'd409,  -13'd254,  -13'd572,  13'd320,  13'd377,  13'd207,  -13'd282,  -13'd94,  -13'd108,  13'd457,  13'd347,  -13'd546,  -13'd416,  
-13'd342,  13'd207,  -13'd296,  -13'd321,  -13'd598,  -13'd170,  13'd301,  -13'd587,  -13'd90,  -13'd214,  -13'd213,  13'd217,  -13'd11,  13'd295,  13'd143,  -13'd678,  
13'd106,  -13'd155,  -13'd331,  -13'd623,  -13'd70,  -13'd236,  13'd630,  13'd58,  13'd746,  13'd118,  -13'd367,  13'd264,  -13'd301,  -13'd213,  -13'd13,  13'd127,  
-13'd6,  13'd214,  -13'd407,  -13'd270,  -13'd255,  13'd446,  13'd87,  13'd454,  13'd185,  13'd137,  13'd304,  13'd215,  13'd65,  -13'd101,  13'd173,  13'd302,  
-13'd142,  -13'd243,  -13'd207,  13'd84,  13'd16,  13'd48,  13'd60,  13'd321,  13'd101,  13'd133,  13'd406,  13'd251,  -13'd691,  -13'd103,  13'd135,  -13'd202,  
13'd306,  -13'd445,  -13'd655,  -13'd837,  -13'd563,  -13'd343,  -13'd235,  -13'd271,  -13'd325,  13'd81,  -13'd160,  -13'd580,  13'd258,  -13'd740,  -13'd374,  -13'd107,  
13'd625,  13'd127,  13'd80,  -13'd166,  13'd152,  -13'd339,  -13'd363,  -13'd125,  -13'd554,  13'd15,  13'd553,  -13'd18,  -13'd388,  -13'd43,  -13'd556,  13'd338,  

13'd355,  13'd148,  -13'd711,  -13'd371,  -13'd1094,  -13'd555,  13'd972,  -13'd1139,  13'd28,  -13'd559,  -13'd735,  -13'd704,  -13'd477,  13'd433,  -13'd943,  -13'd574,  
13'd472,  -13'd123,  13'd628,  -13'd160,  -13'd142,  -13'd192,  13'd145,  13'd351,  -13'd593,  -13'd534,  -13'd721,  -13'd323,  -13'd640,  13'd720,  13'd112,  -13'd1112,  
13'd413,  13'd457,  13'd398,  13'd462,  13'd115,  -13'd636,  13'd276,  13'd329,  13'd177,  13'd134,  13'd562,  13'd144,  13'd212,  -13'd697,  -13'd441,  -13'd1020,  
13'd10,  13'd413,  13'd124,  13'd864,  -13'd1110,  13'd244,  13'd587,  13'd602,  13'd294,  13'd122,  13'd580,  13'd100,  13'd204,  13'd55,  13'd410,  -13'd648,  
-13'd161,  13'd352,  -13'd27,  13'd1023,  -13'd123,  13'd279,  13'd140,  13'd333,  -13'd211,  -13'd193,  13'd311,  -13'd346,  13'd470,  13'd62,  -13'd98,  13'd32,  
-13'd809,  -13'd783,  -13'd554,  -13'd460,  -13'd829,  -13'd874,  13'd223,  -13'd903,  -13'd464,  13'd151,  13'd233,  -13'd532,  -13'd32,  13'd225,  -13'd481,  -13'd729,  
13'd437,  -13'd132,  13'd648,  -13'd427,  -13'd587,  13'd479,  -13'd31,  13'd343,  13'd9,  -13'd149,  -13'd272,  -13'd275,  13'd193,  13'd889,  -13'd76,  -13'd77,  
-13'd448,  -13'd240,  13'd263,  -13'd123,  -13'd27,  13'd314,  13'd284,  13'd894,  13'd753,  13'd488,  13'd361,  -13'd106,  -13'd340,  -13'd1087,  13'd154,  -13'd253,  
-13'd310,  13'd34,  13'd179,  13'd926,  13'd503,  -13'd179,  13'd192,  13'd555,  13'd481,  13'd630,  13'd290,  -13'd704,  13'd837,  13'd50,  -13'd318,  13'd387,  
-13'd828,  -13'd94,  -13'd464,  -13'd238,  -13'd8,  -13'd320,  -13'd1103,  -13'd278,  -13'd647,  13'd388,  13'd692,  13'd258,  13'd293,  -13'd345,  13'd288,  13'd183,  
-13'd27,  -13'd1048,  13'd511,  -13'd230,  -13'd149,  13'd262,  -13'd708,  13'd325,  13'd384,  -13'd479,  -13'd464,  13'd198,  -13'd380,  13'd863,  -13'd145,  -13'd402,  
-13'd42,  -13'd775,  13'd1206,  -13'd465,  -13'd573,  13'd137,  13'd224,  13'd0,  -13'd640,  -13'd82,  13'd153,  -13'd2,  13'd49,  13'd5,  13'd229,  13'd378,  
-13'd491,  -13'd161,  13'd10,  -13'd150,  -13'd271,  13'd90,  13'd144,  13'd46,  -13'd655,  13'd339,  -13'd315,  -13'd420,  13'd443,  -13'd220,  13'd246,  -13'd58,  
-13'd1017,  -13'd527,  13'd1025,  -13'd483,  -13'd87,  -13'd709,  -13'd69,  -13'd66,  -13'd43,  13'd5,  13'd269,  13'd379,  -13'd845,  13'd163,  -13'd2,  -13'd148,  
-13'd1336,  13'd878,  13'd175,  -13'd38,  13'd26,  13'd263,  -13'd40,  -13'd16,  13'd32,  -13'd127,  13'd578,  -13'd389,  -13'd1418,  -13'd317,  -13'd345,  -13'd600,  
-13'd199,  13'd195,  -13'd632,  -13'd137,  13'd776,  13'd241,  -13'd1374,  -13'd405,  -13'd277,  13'd109,  -13'd387,  -13'd493,  -13'd340,  13'd7,  -13'd28,  -13'd503,  
13'd77,  -13'd465,  13'd300,  13'd516,  13'd318,  -13'd245,  -13'd352,  -13'd180,  -13'd1294,  -13'd105,  -13'd841,  13'd279,  -13'd168,  13'd266,  13'd58,  13'd163,  
13'd437,  13'd173,  13'd452,  -13'd64,  -13'd347,  13'd94,  13'd655,  -13'd11,  -13'd142,  -13'd454,  -13'd580,  -13'd122,  13'd207,  13'd721,  13'd439,  -13'd67,  
-13'd710,  -13'd389,  13'd818,  13'd518,  -13'd86,  -13'd318,  13'd604,  13'd828,  13'd293,  -13'd428,  -13'd38,  -13'd328,  -13'd277,  -13'd372,  -13'd364,  -13'd175,  
-13'd95,  13'd253,  13'd1099,  -13'd866,  -13'd266,  -13'd197,  -13'd395,  13'd298,  -13'd68,  -13'd528,  -13'd181,  -13'd643,  -13'd250,  13'd288,  -13'd549,  -13'd716,  
-13'd916,  13'd109,  -13'd628,  13'd753,  13'd128,  13'd110,  13'd114,  13'd426,  13'd658,  13'd122,  13'd524,  -13'd225,  13'd188,  -13'd1027,  13'd57,  -13'd203,  
13'd226,  -13'd235,  13'd39,  13'd461,  13'd439,  -13'd154,  -13'd357,  -13'd390,  13'd660,  13'd2,  13'd847,  -13'd108,  13'd206,  -13'd978,  -13'd63,  -13'd72,  
13'd488,  13'd495,  13'd539,  -13'd12,  13'd377,  13'd91,  -13'd341,  13'd48,  -13'd292,  13'd656,  13'd53,  13'd136,  -13'd682,  13'd712,  13'd217,  -13'd157,  
-13'd799,  13'd19,  13'd112,  13'd651,  -13'd544,  -13'd356,  13'd639,  -13'd121,  -13'd381,  -13'd578,  13'd351,  -13'd358,  -13'd251,  -13'd641,  13'd57,  -13'd238,  
-13'd486,  -13'd930,  -13'd837,  -13'd380,  -13'd860,  -13'd1319,  13'd410,  -13'd578,  13'd352,  -13'd90,  -13'd651,  -13'd158,  -13'd324,  13'd382,  -13'd225,  -13'd806,  

13'd39,  13'd230,  13'd634,  13'd469,  -13'd334,  -13'd804,  13'd315,  -13'd84,  -13'd254,  -13'd35,  13'd528,  -13'd593,  -13'd307,  -13'd5,  -13'd629,  -13'd129,  
13'd352,  -13'd127,  -13'd100,  -13'd131,  -13'd786,  13'd470,  13'd183,  -13'd359,  -13'd222,  -13'd621,  13'd278,  -13'd407,  -13'd142,  -13'd619,  -13'd665,  13'd287,  
-13'd194,  13'd285,  13'd99,  13'd311,  -13'd629,  -13'd437,  -13'd45,  -13'd427,  13'd23,  -13'd350,  13'd227,  13'd343,  -13'd110,  13'd249,  13'd156,  13'd10,  
-13'd287,  13'd404,  -13'd520,  13'd28,  13'd460,  -13'd882,  13'd209,  -13'd33,  -13'd338,  -13'd565,  13'd563,  13'd101,  13'd0,  -13'd230,  13'd311,  13'd52,  
13'd302,  13'd346,  -13'd391,  -13'd46,  13'd530,  -13'd155,  -13'd278,  -13'd104,  13'd148,  13'd239,  13'd608,  -13'd461,  -13'd25,  13'd429,  -13'd447,  13'd462,  
-13'd584,  -13'd371,  13'd195,  -13'd56,  -13'd423,  -13'd319,  13'd256,  -13'd107,  -13'd136,  13'd371,  13'd298,  -13'd381,  -13'd370,  13'd239,  -13'd257,  13'd16,  
13'd277,  -13'd257,  -13'd24,  -13'd454,  -13'd435,  -13'd57,  -13'd366,  -13'd359,  -13'd187,  -13'd55,  13'd576,  -13'd269,  -13'd425,  13'd225,  13'd69,  -13'd311,  
-13'd161,  13'd166,  -13'd313,  -13'd486,  13'd394,  -13'd168,  -13'd289,  -13'd484,  -13'd73,  13'd24,  -13'd127,  13'd302,  -13'd391,  13'd698,  -13'd808,  -13'd756,  
-13'd646,  13'd259,  -13'd575,  13'd176,  -13'd124,  -13'd345,  -13'd376,  13'd323,  -13'd323,  -13'd599,  -13'd862,  -13'd62,  -13'd15,  13'd112,  -13'd13,  13'd96,  
13'd113,  13'd552,  -13'd246,  13'd313,  -13'd523,  -13'd173,  -13'd4,  -13'd542,  13'd581,  -13'd152,  13'd75,  -13'd633,  -13'd73,  13'd153,  13'd474,  -13'd321,  
-13'd585,  13'd156,  13'd290,  -13'd647,  13'd73,  -13'd65,  -13'd625,  13'd326,  -13'd126,  13'd164,  -13'd369,  -13'd282,  13'd108,  -13'd591,  -13'd332,  -13'd8,  
-13'd463,  -13'd807,  -13'd11,  -13'd169,  -13'd816,  -13'd624,  -13'd290,  -13'd695,  -13'd311,  -13'd278,  -13'd45,  13'd392,  13'd81,  -13'd68,  -13'd155,  13'd265,  
-13'd225,  -13'd218,  13'd443,  -13'd395,  -13'd647,  -13'd578,  13'd193,  -13'd62,  -13'd23,  -13'd329,  -13'd488,  -13'd805,  -13'd73,  -13'd85,  -13'd292,  -13'd154,  
13'd40,  13'd332,  -13'd497,  13'd580,  -13'd462,  -13'd120,  -13'd519,  -13'd290,  13'd224,  -13'd14,  -13'd194,  -13'd308,  13'd210,  13'd242,  -13'd54,  13'd344,  
-13'd218,  13'd209,  -13'd30,  -13'd225,  13'd8,  13'd58,  -13'd229,  13'd234,  -13'd488,  -13'd176,  -13'd728,  -13'd726,  13'd153,  13'd510,  13'd67,  13'd215,  
-13'd211,  13'd41,  -13'd109,  13'd535,  13'd431,  -13'd36,  -13'd178,  -13'd368,  13'd166,  -13'd326,  13'd501,  13'd520,  -13'd114,  -13'd207,  -13'd501,  13'd336,  
13'd168,  -13'd18,  -13'd455,  -13'd2,  13'd27,  -13'd644,  -13'd36,  13'd208,  13'd210,  -13'd158,  -13'd471,  -13'd318,  -13'd476,  -13'd112,  -13'd322,  13'd297,  
13'd284,  -13'd21,  -13'd456,  13'd427,  13'd105,  13'd156,  13'd90,  13'd43,  -13'd180,  13'd594,  13'd720,  -13'd719,  -13'd113,  -13'd49,  -13'd470,  13'd31,  
-13'd202,  -13'd164,  -13'd178,  -13'd483,  -13'd553,  -13'd405,  -13'd457,  -13'd80,  -13'd602,  13'd118,  13'd349,  -13'd816,  13'd408,  -13'd825,  13'd110,  -13'd423,  
13'd742,  -13'd194,  13'd238,  -13'd246,  13'd219,  -13'd650,  -13'd582,  -13'd704,  -13'd247,  13'd190,  13'd381,  13'd558,  -13'd433,  13'd16,  -13'd303,  13'd65,  
-13'd82,  13'd76,  13'd198,  -13'd84,  13'd55,  13'd662,  -13'd141,  13'd19,  -13'd141,  -13'd628,  13'd314,  -13'd239,  13'd81,  13'd285,  13'd102,  -13'd184,  
-13'd680,  -13'd294,  -13'd293,  -13'd150,  13'd232,  13'd100,  -13'd4,  13'd103,  -13'd507,  -13'd471,  13'd287,  13'd179,  13'd560,  13'd330,  -13'd794,  13'd253,  
-13'd235,  -13'd95,  13'd357,  -13'd847,  -13'd567,  -13'd848,  -13'd41,  13'd479,  -13'd336,  -13'd463,  13'd106,  13'd132,  -13'd322,  -13'd162,  13'd631,  13'd69,  
-13'd39,  -13'd492,  13'd535,  -13'd107,  -13'd608,  -13'd343,  13'd135,  13'd93,  -13'd3,  -13'd101,  -13'd588,  -13'd301,  13'd496,  13'd111,  13'd82,  13'd254,  
-13'd175,  -13'd514,  13'd168,  13'd356,  -13'd14,  13'd56,  -13'd25,  13'd71,  -13'd133,  -13'd218,  -13'd279,  13'd140,  13'd288,  -13'd385,  13'd258,  13'd204,  

-13'd206,  -13'd786,  13'd70,  13'd79,  -13'd64,  -13'd323,  13'd570,  13'd783,  13'd413,  13'd157,  13'd296,  -13'd846,  13'd341,  -13'd350,  13'd395,  13'd154,  
13'd513,  13'd161,  -13'd5,  -13'd609,  13'd573,  -13'd45,  -13'd88,  13'd823,  -13'd151,  13'd597,  13'd503,  -13'd56,  13'd850,  -13'd556,  13'd398,  -13'd748,  
13'd6,  -13'd610,  13'd125,  13'd457,  -13'd537,  13'd280,  13'd2,  -13'd140,  13'd0,  13'd20,  -13'd132,  13'd307,  13'd665,  -13'd404,  13'd23,  -13'd90,  
13'd920,  -13'd25,  13'd597,  -13'd72,  -13'd377,  -13'd556,  13'd233,  13'd133,  13'd660,  -13'd593,  13'd28,  -13'd341,  13'd980,  -13'd475,  13'd809,  -13'd75,  
-13'd268,  -13'd455,  13'd261,  -13'd606,  -13'd173,  -13'd419,  -13'd530,  13'd648,  13'd55,  -13'd100,  13'd431,  13'd412,  13'd411,  -13'd415,  -13'd369,  13'd6,  
-13'd58,  13'd412,  13'd340,  13'd558,  13'd747,  -13'd355,  -13'd855,  -13'd315,  -13'd113,  -13'd76,  -13'd119,  13'd73,  -13'd95,  -13'd34,  -13'd707,  -13'd104,  
-13'd716,  13'd877,  13'd64,  -13'd297,  -13'd326,  13'd516,  -13'd509,  -13'd505,  13'd551,  -13'd56,  -13'd155,  -13'd172,  13'd7,  -13'd6,  -13'd481,  -13'd407,  
-13'd732,  13'd822,  -13'd205,  13'd232,  13'd460,  13'd369,  13'd79,  -13'd0,  -13'd234,  13'd200,  13'd481,  -13'd201,  13'd385,  13'd189,  13'd264,  13'd781,  
-13'd343,  13'd728,  -13'd49,  13'd26,  13'd256,  -13'd434,  -13'd587,  -13'd53,  13'd170,  -13'd396,  13'd289,  -13'd66,  13'd454,  13'd145,  13'd308,  13'd169,  
-13'd387,  13'd222,  13'd171,  13'd335,  -13'd498,  13'd258,  -13'd703,  -13'd483,  -13'd114,  13'd330,  -13'd451,  13'd1073,  13'd535,  -13'd240,  13'd302,  13'd691,  
-13'd169,  13'd126,  13'd14,  -13'd504,  -13'd7,  -13'd83,  -13'd544,  13'd41,  13'd460,  -13'd504,  13'd1131,  13'd448,  13'd164,  13'd24,  13'd388,  -13'd529,  
13'd543,  13'd436,  13'd891,  -13'd632,  -13'd249,  -13'd398,  -13'd60,  -13'd652,  13'd397,  13'd74,  13'd70,  -13'd50,  -13'd528,  -13'd34,  -13'd543,  13'd431,  
13'd191,  13'd118,  -13'd268,  13'd5,  -13'd110,  -13'd227,  13'd101,  -13'd127,  -13'd339,  -13'd188,  13'd16,  -13'd551,  13'd111,  13'd279,  13'd90,  13'd8,  
-13'd451,  13'd339,  -13'd422,  -13'd406,  13'd954,  13'd468,  13'd56,  -13'd544,  -13'd386,  13'd169,  13'd151,  13'd382,  13'd444,  -13'd30,  -13'd45,  13'd62,  
13'd71,  13'd244,  13'd1388,  13'd257,  13'd821,  -13'd854,  13'd223,  13'd48,  13'd321,  13'd712,  13'd419,  13'd588,  -13'd380,  13'd16,  13'd53,  13'd682,  
13'd647,  13'd206,  13'd203,  -13'd479,  -13'd139,  -13'd692,  13'd348,  13'd22,  -13'd141,  -13'd466,  13'd454,  -13'd198,  -13'd573,  13'd83,  13'd84,  13'd1,  
13'd615,  13'd88,  13'd43,  13'd48,  13'd202,  -13'd449,  13'd469,  -13'd262,  13'd203,  13'd302,  -13'd315,  13'd235,  13'd310,  13'd586,  -13'd364,  -13'd148,  
-13'd175,  -13'd143,  13'd264,  -13'd654,  -13'd255,  13'd441,  13'd351,  13'd135,  13'd319,  -13'd700,  -13'd89,  13'd752,  13'd48,  -13'd345,  -13'd296,  -13'd443,  
-13'd100,  -13'd475,  13'd4,  -13'd121,  -13'd457,  13'd373,  13'd468,  -13'd212,  -13'd211,  -13'd227,  -13'd282,  13'd251,  13'd207,  13'd190,  -13'd827,  13'd28,  
-13'd260,  13'd50,  13'd745,  13'd284,  -13'd773,  13'd171,  13'd491,  13'd414,  13'd288,  -13'd370,  -13'd190,  -13'd223,  13'd583,  -13'd227,  13'd401,  -13'd538,  
-13'd214,  -13'd41,  13'd181,  13'd268,  -13'd306,  -13'd153,  -13'd48,  13'd518,  -13'd175,  -13'd69,  -13'd524,  -13'd606,  13'd202,  13'd629,  -13'd213,  13'd555,  
13'd140,  -13'd15,  13'd382,  13'd334,  -13'd425,  13'd348,  -13'd605,  13'd629,  -13'd536,  13'd580,  13'd119,  13'd400,  13'd221,  13'd248,  13'd908,  -13'd99,  
13'd589,  13'd158,  -13'd262,  13'd59,  13'd158,  13'd326,  -13'd311,  -13'd498,  13'd381,  -13'd302,  13'd580,  13'd210,  13'd121,  -13'd98,  -13'd517,  -13'd197,  
13'd118,  -13'd214,  13'd344,  -13'd716,  13'd147,  -13'd238,  13'd559,  -13'd341,  -13'd437,  13'd54,  -13'd31,  13'd283,  -13'd264,  13'd231,  -13'd97,  13'd264,  
13'd387,  13'd210,  13'd805,  -13'd587,  -13'd597,  -13'd94,  13'd3,  -13'd109,  13'd87,  -13'd101,  -13'd501,  -13'd281,  -13'd868,  13'd660,  -13'd409,  -13'd289,  

13'd102,  13'd518,  13'd264,  -13'd123,  13'd190,  13'd137,  13'd538,  13'd263,  -13'd177,  -13'd24,  13'd202,  -13'd3,  13'd314,  13'd332,  13'd704,  -13'd6,  
13'd1049,  13'd217,  13'd837,  -13'd226,  -13'd484,  13'd237,  13'd745,  -13'd378,  -13'd14,  -13'd616,  13'd503,  13'd369,  -13'd41,  13'd794,  -13'd234,  13'd573,  
13'd289,  -13'd214,  13'd695,  -13'd397,  -13'd574,  -13'd434,  13'd1034,  -13'd739,  -13'd852,  -13'd429,  13'd309,  -13'd748,  13'd130,  13'd160,  -13'd722,  -13'd356,  
-13'd388,  -13'd22,  -13'd1344,  -13'd1027,  -13'd82,  -13'd678,  13'd946,  -13'd733,  -13'd524,  -13'd1127,  13'd886,  -13'd22,  -13'd161,  13'd587,  -13'd418,  -13'd86,  
-13'd489,  13'd145,  -13'd1101,  -13'd593,  -13'd679,  -13'd440,  -13'd1137,  -13'd1099,  -13'd987,  -13'd278,  -13'd60,  -13'd704,  -13'd1040,  -13'd161,  -13'd550,  13'd467,  
13'd854,  -13'd61,  13'd289,  -13'd6,  -13'd409,  -13'd477,  13'd29,  13'd33,  13'd723,  -13'd600,  13'd682,  13'd653,  13'd997,  13'd52,  13'd444,  13'd129,  
-13'd31,  13'd568,  -13'd221,  -13'd602,  13'd415,  -13'd553,  13'd423,  13'd9,  -13'd520,  13'd611,  13'd477,  -13'd302,  -13'd70,  13'd273,  13'd79,  13'd73,  
-13'd156,  -13'd798,  13'd289,  -13'd305,  -13'd309,  -13'd1465,  -13'd99,  -13'd576,  13'd175,  -13'd36,  13'd110,  13'd354,  -13'd178,  -13'd523,  -13'd709,  -13'd709,  
13'd174,  13'd168,  -13'd566,  -13'd92,  -13'd564,  13'd126,  -13'd314,  -13'd1094,  13'd827,  13'd713,  -13'd389,  -13'd474,  -13'd302,  -13'd361,  -13'd618,  -13'd683,  
13'd836,  -13'd904,  -13'd12,  13'd502,  13'd627,  -13'd213,  -13'd6,  -13'd902,  13'd238,  13'd686,  -13'd674,  13'd885,  13'd90,  13'd34,  -13'd396,  13'd78,  
-13'd383,  13'd27,  13'd672,  13'd139,  -13'd450,  -13'd500,  13'd374,  -13'd111,  -13'd231,  13'd35,  -13'd4,  -13'd298,  -13'd648,  13'd10,  -13'd535,  13'd328,  
-13'd613,  13'd716,  13'd876,  -13'd609,  -13'd289,  -13'd379,  13'd135,  -13'd148,  13'd224,  -13'd347,  -13'd474,  -13'd725,  -13'd707,  13'd627,  13'd125,  -13'd1089,  
13'd475,  -13'd1198,  13'd423,  13'd92,  -13'd667,  -13'd457,  -13'd689,  -13'd481,  -13'd531,  13'd193,  -13'd489,  -13'd53,  -13'd1217,  -13'd32,  -13'd297,  13'd181,  
13'd825,  -13'd283,  -13'd1057,  13'd268,  13'd36,  13'd488,  -13'd489,  -13'd102,  13'd888,  13'd153,  13'd913,  13'd422,  13'd366,  -13'd19,  -13'd127,  13'd557,  
13'd560,  13'd319,  13'd156,  13'd254,  13'd700,  13'd652,  13'd473,  -13'd110,  13'd517,  13'd507,  13'd1106,  13'd578,  13'd374,  -13'd102,  13'd478,  13'd343,  
-13'd414,  13'd216,  -13'd586,  -13'd4,  13'd504,  -13'd309,  13'd180,  13'd297,  13'd346,  -13'd840,  -13'd366,  -13'd413,  13'd424,  -13'd187,  13'd227,  13'd265,  
13'd58,  -13'd381,  13'd317,  13'd264,  -13'd308,  13'd555,  -13'd256,  13'd328,  -13'd317,  -13'd105,  13'd423,  -13'd127,  13'd65,  13'd649,  13'd26,  -13'd380,  
13'd274,  -13'd763,  13'd604,  13'd534,  -13'd160,  -13'd180,  -13'd219,  13'd518,  -13'd1065,  13'd181,  13'd464,  -13'd85,  13'd805,  -13'd281,  13'd392,  -13'd1017,  
-13'd36,  -13'd281,  -13'd505,  13'd768,  13'd733,  -13'd15,  13'd551,  13'd470,  -13'd860,  -13'd300,  13'd615,  13'd409,  13'd358,  -13'd418,  13'd739,  -13'd27,  
-13'd111,  13'd68,  -13'd270,  13'd410,  -13'd254,  13'd99,  13'd353,  13'd876,  -13'd373,  13'd618,  13'd383,  13'd148,  13'd904,  -13'd136,  13'd112,  13'd388,  
13'd98,  -13'd99,  13'd75,  13'd24,  13'd467,  -13'd328,  -13'd937,  13'd263,  13'd141,  13'd98,  13'd33,  -13'd1031,  13'd245,  -13'd50,  -13'd674,  -13'd280,  
-13'd865,  13'd407,  -13'd293,  13'd366,  -13'd264,  -13'd57,  -13'd1384,  13'd254,  13'd750,  13'd166,  13'd316,  -13'd1182,  13'd510,  13'd458,  -13'd524,  13'd241,  
13'd19,  -13'd354,  -13'd1206,  13'd95,  -13'd458,  13'd486,  -13'd222,  13'd142,  -13'd1022,  -13'd226,  13'd655,  13'd10,  13'd601,  -13'd1805,  -13'd547,  -13'd421,  
-13'd838,  -13'd762,  -13'd2010,  13'd65,  13'd403,  -13'd193,  -13'd233,  -13'd55,  13'd290,  -13'd936,  13'd494,  13'd15,  13'd69,  -13'd84,  -13'd796,  13'd2,  
13'd77,  -13'd833,  -13'd677,  -13'd728,  13'd174,  -13'd1057,  -13'd689,  13'd468,  -13'd148,  13'd1017,  13'd18,  -13'd636,  -13'd603,  -13'd473,  -13'd454,  13'd369,  

-13'd338,  -13'd293,  13'd658,  13'd454,  -13'd124,  -13'd258,  -13'd591,  13'd183,  13'd139,  -13'd197,  -13'd303,  -13'd243,  -13'd329,  -13'd316,  13'd324,  -13'd173,  
13'd758,  -13'd462,  13'd314,  13'd807,  13'd224,  13'd858,  -13'd165,  13'd239,  -13'd445,  -13'd471,  -13'd597,  13'd59,  13'd713,  13'd293,  13'd504,  -13'd1089,  
-13'd330,  13'd199,  -13'd184,  -13'd273,  -13'd225,  13'd919,  -13'd320,  13'd607,  13'd1192,  13'd590,  -13'd32,  -13'd610,  13'd542,  -13'd512,  13'd830,  -13'd577,  
-13'd79,  -13'd232,  -13'd477,  13'd113,  -13'd420,  -13'd418,  -13'd1006,  -13'd30,  -13'd863,  13'd375,  -13'd483,  -13'd648,  13'd2,  -13'd687,  13'd243,  13'd787,  
-13'd60,  -13'd399,  13'd355,  13'd85,  13'd280,  -13'd95,  13'd294,  13'd630,  -13'd47,  13'd282,  -13'd42,  13'd250,  13'd26,  -13'd406,  -13'd109,  -13'd654,  
13'd492,  -13'd80,  13'd119,  -13'd383,  -13'd597,  13'd184,  13'd80,  -13'd256,  -13'd216,  13'd93,  -13'd65,  13'd398,  -13'd220,  13'd645,  13'd488,  -13'd398,  
13'd318,  -13'd532,  13'd1370,  13'd279,  -13'd77,  13'd728,  -13'd368,  13'd128,  13'd503,  -13'd768,  -13'd670,  -13'd658,  -13'd126,  13'd37,  -13'd679,  -13'd417,  
-13'd414,  13'd1010,  -13'd708,  -13'd422,  13'd260,  13'd1161,  -13'd192,  13'd780,  13'd870,  -13'd300,  -13'd10,  13'd104,  13'd313,  13'd343,  13'd42,  13'd275,  
13'd251,  13'd325,  -13'd196,  13'd152,  13'd142,  13'd272,  -13'd599,  13'd547,  -13'd578,  -13'd55,  -13'd254,  -13'd603,  13'd441,  13'd249,  13'd721,  -13'd359,  
-13'd87,  -13'd438,  13'd72,  13'd153,  13'd651,  13'd133,  13'd24,  13'd209,  -13'd454,  13'd371,  13'd723,  13'd1157,  13'd115,  -13'd589,  13'd102,  13'd488,  
13'd389,  -13'd292,  13'd719,  13'd472,  13'd115,  13'd727,  -13'd48,  13'd134,  -13'd229,  -13'd172,  -13'd35,  13'd370,  -13'd559,  13'd117,  -13'd444,  -13'd455,  
13'd379,  13'd991,  -13'd22,  -13'd245,  13'd288,  13'd460,  13'd523,  -13'd441,  -13'd4,  -13'd618,  13'd90,  13'd163,  13'd520,  -13'd435,  -13'd514,  -13'd132,  
13'd269,  13'd772,  -13'd751,  13'd117,  13'd641,  -13'd51,  13'd495,  -13'd631,  -13'd435,  -13'd140,  -13'd671,  -13'd1007,  -13'd539,  13'd399,  13'd99,  -13'd546,  
13'd417,  13'd897,  -13'd446,  -13'd948,  13'd467,  13'd7,  -13'd377,  13'd28,  -13'd203,  -13'd448,  -13'd418,  13'd110,  -13'd106,  13'd276,  13'd753,  13'd271,  
13'd211,  13'd634,  13'd133,  -13'd79,  13'd575,  -13'd176,  -13'd35,  -13'd177,  -13'd369,  -13'd1697,  13'd386,  -13'd352,  13'd4,  -13'd480,  13'd273,  13'd28,  
13'd385,  -13'd291,  13'd256,  13'd620,  13'd72,  -13'd195,  13'd100,  13'd576,  -13'd485,  -13'd280,  -13'd552,  -13'd65,  -13'd508,  -13'd211,  13'd328,  -13'd127,  
13'd18,  -13'd211,  -13'd186,  -13'd573,  -13'd173,  -13'd251,  13'd1173,  13'd593,  -13'd98,  -13'd833,  -13'd423,  -13'd234,  -13'd846,  13'd95,  13'd494,  -13'd808,  
13'd503,  13'd314,  13'd422,  13'd244,  -13'd142,  -13'd312,  -13'd162,  -13'd119,  13'd442,  13'd50,  -13'd24,  -13'd78,  -13'd444,  13'd740,  -13'd65,  -13'd619,  
13'd543,  13'd541,  13'd191,  -13'd202,  13'd24,  13'd493,  13'd353,  -13'd104,  13'd10,  13'd262,  13'd217,  13'd535,  13'd270,  13'd716,  -13'd676,  -13'd279,  
13'd413,  13'd397,  13'd534,  -13'd331,  13'd150,  13'd524,  13'd517,  13'd427,  -13'd159,  -13'd218,  13'd115,  13'd223,  -13'd77,  -13'd86,  -13'd1009,  13'd256,  
-13'd519,  13'd530,  13'd125,  13'd1,  -13'd702,  13'd289,  -13'd186,  13'd569,  13'd110,  -13'd117,  -13'd143,  13'd568,  -13'd417,  -13'd367,  -13'd427,  13'd98,  
13'd165,  -13'd159,  -13'd379,  -13'd139,  13'd68,  13'd452,  13'd131,  13'd69,  13'd132,  13'd212,  13'd7,  13'd218,  13'd408,  -13'd300,  13'd110,  -13'd139,  
-13'd298,  -13'd742,  -13'd354,  -13'd211,  13'd199,  13'd114,  -13'd284,  -13'd102,  13'd238,  13'd90,  -13'd260,  13'd435,  -13'd51,  -13'd302,  -13'd645,  13'd108,  
13'd1239,  -13'd740,  13'd869,  -13'd220,  13'd439,  13'd16,  -13'd370,  13'd258,  13'd353,  13'd272,  13'd469,  13'd581,  13'd215,  -13'd227,  -13'd1181,  -13'd468,  
13'd1004,  13'd487,  -13'd217,  -13'd967,  -13'd219,  -13'd689,  -13'd494,  13'd92,  -13'd540,  -13'd818,  -13'd877,  -13'd440,  13'd126,  -13'd331,  -13'd1119,  13'd257,  

13'd751,  13'd306,  -13'd595,  -13'd25,  -13'd225,  -13'd336,  13'd455,  -13'd341,  13'd590,  -13'd311,  -13'd355,  13'd164,  -13'd1025,  -13'd297,  13'd273,  -13'd677,  
13'd522,  13'd300,  13'd95,  -13'd351,  -13'd431,  13'd7,  -13'd171,  13'd450,  -13'd250,  13'd627,  -13'd241,  -13'd341,  -13'd113,  -13'd114,  13'd137,  -13'd176,  
13'd383,  -13'd303,  -13'd180,  13'd45,  13'd15,  13'd112,  -13'd771,  -13'd529,  13'd2,  13'd851,  -13'd68,  13'd43,  -13'd567,  -13'd206,  13'd202,  13'd693,  
-13'd229,  -13'd455,  13'd285,  13'd346,  -13'd284,  -13'd453,  -13'd192,  -13'd328,  13'd283,  13'd151,  13'd515,  -13'd856,  13'd549,  -13'd631,  -13'd123,  13'd48,  
13'd606,  -13'd392,  13'd109,  -13'd28,  13'd797,  -13'd274,  -13'd324,  13'd407,  -13'd437,  -13'd327,  13'd237,  13'd189,  -13'd292,  13'd84,  -13'd18,  13'd1149,  
13'd118,  -13'd144,  13'd539,  -13'd163,  13'd646,  13'd314,  -13'd508,  -13'd41,  13'd422,  13'd827,  -13'd468,  -13'd40,  -13'd223,  -13'd369,  13'd981,  13'd111,  
-13'd305,  13'd495,  13'd319,  13'd36,  13'd222,  -13'd248,  -13'd141,  13'd831,  13'd107,  13'd372,  -13'd828,  -13'd472,  13'd212,  13'd340,  13'd781,  13'd1048,  
-13'd213,  -13'd12,  13'd115,  13'd557,  -13'd733,  -13'd77,  -13'd356,  13'd268,  13'd143,  -13'd471,  13'd174,  -13'd29,  13'd455,  -13'd592,  -13'd337,  13'd56,  
-13'd498,  -13'd354,  -13'd497,  -13'd26,  -13'd412,  -13'd164,  13'd96,  13'd122,  -13'd145,  13'd123,  -13'd318,  13'd560,  -13'd300,  -13'd979,  -13'd355,  13'd273,  
-13'd16,  13'd756,  -13'd440,  -13'd252,  -13'd0,  13'd377,  -13'd33,  13'd782,  -13'd291,  13'd360,  -13'd308,  13'd334,  13'd908,  13'd44,  -13'd550,  13'd9,  
-13'd267,  -13'd368,  -13'd426,  13'd846,  13'd926,  13'd178,  -13'd1857,  13'd634,  -13'd2,  13'd911,  13'd33,  13'd975,  -13'd194,  -13'd295,  -13'd63,  13'd47,  
-13'd211,  13'd1235,  13'd474,  13'd123,  -13'd29,  13'd522,  -13'd406,  13'd100,  -13'd149,  13'd782,  13'd882,  13'd518,  -13'd13,  13'd113,  -13'd69,  13'd574,  
13'd219,  13'd30,  -13'd3,  13'd424,  -13'd374,  13'd5,  -13'd635,  -13'd288,  -13'd93,  13'd157,  13'd520,  13'd706,  13'd13,  -13'd528,  -13'd146,  13'd185,  
-13'd586,  -13'd443,  13'd32,  -13'd422,  13'd655,  -13'd816,  13'd385,  13'd197,  -13'd290,  -13'd57,  13'd372,  13'd178,  13'd472,  13'd375,  -13'd50,  13'd768,  
13'd782,  -13'd276,  -13'd706,  -13'd81,  13'd141,  13'd8,  -13'd275,  -13'd710,  -13'd309,  -13'd11,  -13'd68,  -13'd295,  13'd261,  -13'd176,  -13'd214,  13'd403,  
-13'd70,  -13'd649,  -13'd148,  13'd412,  13'd1373,  -13'd51,  -13'd702,  13'd251,  13'd292,  13'd469,  -13'd220,  13'd836,  -13'd174,  13'd423,  13'd491,  13'd70,  
13'd492,  13'd270,  -13'd213,  13'd350,  13'd681,  -13'd16,  13'd135,  -13'd852,  13'd861,  13'd981,  -13'd372,  13'd469,  13'd712,  -13'd48,  -13'd132,  13'd287,  
-13'd217,  13'd716,  13'd70,  -13'd265,  13'd167,  -13'd822,  13'd345,  -13'd136,  13'd724,  -13'd336,  -13'd369,  13'd257,  -13'd625,  13'd372,  -13'd322,  -13'd556,  
13'd219,  -13'd83,  13'd72,  -13'd737,  13'd10,  -13'd10,  -13'd569,  -13'd302,  -13'd91,  -13'd172,  -13'd1072,  13'd123,  13'd180,  13'd86,  -13'd316,  -13'd786,  
-13'd350,  -13'd78,  13'd878,  -13'd22,  -13'd154,  13'd134,  13'd141,  -13'd168,  13'd203,  13'd75,  -13'd809,  13'd427,  -13'd328,  13'd23,  13'd393,  -13'd799,  
13'd250,  13'd168,  -13'd12,  -13'd78,  13'd134,  13'd770,  13'd593,  13'd987,  13'd337,  -13'd50,  -13'd53,  13'd630,  13'd113,  13'd124,  13'd32,  13'd474,  
-13'd72,  -13'd116,  -13'd546,  13'd276,  -13'd30,  -13'd74,  -13'd1001,  13'd622,  -13'd604,  -13'd8,  -13'd103,  -13'd524,  13'd301,  13'd351,  13'd523,  -13'd160,  
13'd433,  -13'd776,  -13'd306,  -13'd192,  -13'd576,  -13'd388,  13'd306,  -13'd164,  13'd115,  13'd787,  13'd57,  13'd929,  13'd216,  -13'd29,  13'd280,  -13'd371,  
13'd92,  -13'd247,  -13'd196,  13'd584,  -13'd353,  13'd719,  -13'd628,  -13'd659,  13'd261,  -13'd29,  13'd558,  13'd629,  -13'd1,  13'd301,  13'd105,  -13'd183,  
13'd788,  -13'd264,  13'd1347,  13'd651,  -13'd314,  13'd996,  -13'd84,  13'd289,  13'd798,  -13'd238,  -13'd115,  13'd266,  -13'd119,  13'd7,  13'd826,  -13'd482,  

-13'd261,  13'd366,  -13'd251,  -13'd348,  -13'd102,  13'd192,  13'd194,  13'd594,  13'd470,  -13'd69,  13'd28,  -13'd131,  13'd1104,  13'd399,  13'd95,  -13'd174,  
13'd451,  13'd589,  13'd913,  -13'd35,  13'd64,  13'd235,  13'd249,  13'd107,  13'd243,  13'd20,  13'd260,  -13'd614,  13'd350,  13'd177,  13'd255,  13'd431,  
-13'd314,  -13'd363,  13'd207,  13'd321,  -13'd65,  13'd72,  13'd314,  13'd445,  13'd131,  13'd34,  -13'd152,  13'd185,  13'd261,  -13'd207,  -13'd286,  13'd483,  
13'd384,  13'd93,  13'd632,  13'd243,  -13'd522,  13'd299,  -13'd463,  -13'd44,  -13'd240,  -13'd168,  -13'd358,  13'd234,  13'd489,  -13'd351,  -13'd78,  13'd61,  
13'd211,  13'd395,  13'd140,  -13'd196,  -13'd278,  -13'd38,  13'd122,  -13'd9,  -13'd159,  -13'd422,  -13'd401,  13'd500,  -13'd213,  -13'd335,  13'd276,  -13'd627,  
-13'd474,  13'd194,  -13'd336,  13'd275,  13'd38,  13'd149,  -13'd378,  -13'd720,  -13'd179,  -13'd747,  13'd513,  13'd332,  13'd7,  13'd629,  -13'd1,  13'd465,  
-13'd217,  13'd8,  13'd891,  -13'd409,  -13'd370,  13'd691,  13'd510,  -13'd937,  -13'd8,  -13'd293,  13'd733,  13'd57,  13'd79,  13'd346,  -13'd616,  13'd169,  
13'd23,  13'd1127,  -13'd564,  13'd418,  13'd271,  13'd766,  13'd1110,  -13'd472,  13'd87,  13'd169,  13'd66,  -13'd51,  -13'd180,  13'd433,  -13'd130,  13'd786,  
13'd2,  13'd689,  13'd107,  -13'd549,  13'd890,  -13'd200,  -13'd301,  13'd262,  -13'd439,  13'd459,  -13'd57,  13'd55,  13'd624,  -13'd338,  13'd212,  13'd98,  
13'd1194,  13'd249,  -13'd318,  -13'd783,  -13'd302,  -13'd425,  -13'd77,  -13'd400,  13'd648,  13'd930,  13'd132,  13'd498,  -13'd166,  -13'd520,  13'd229,  13'd31,  
-13'd175,  -13'd356,  -13'd165,  -13'd388,  -13'd780,  -13'd444,  13'd393,  13'd459,  -13'd302,  -13'd81,  13'd286,  13'd340,  13'd372,  -13'd240,  13'd87,  -13'd157,  
13'd607,  13'd225,  13'd38,  -13'd371,  13'd33,  -13'd536,  13'd373,  -13'd344,  -13'd548,  -13'd563,  -13'd225,  -13'd246,  13'd24,  13'd73,  13'd128,  -13'd37,  
-13'd16,  13'd1186,  13'd329,  -13'd692,  13'd298,  -13'd642,  13'd574,  -13'd41,  -13'd136,  13'd374,  -13'd786,  -13'd203,  -13'd1251,  13'd1218,  -13'd7,  13'd512,  
-13'd296,  13'd590,  13'd491,  -13'd185,  13'd53,  -13'd197,  13'd185,  13'd416,  13'd38,  -13'd567,  13'd71,  13'd58,  -13'd1105,  13'd476,  13'd139,  -13'd735,  
13'd82,  13'd86,  13'd506,  -13'd875,  -13'd786,  -13'd43,  13'd513,  -13'd25,  -13'd175,  -13'd506,  -13'd450,  -13'd216,  -13'd463,  -13'd463,  13'd1030,  -13'd742,  
13'd1137,  13'd89,  13'd124,  -13'd1181,  -13'd516,  -13'd387,  13'd38,  -13'd725,  -13'd474,  13'd27,  -13'd784,  13'd541,  -13'd1331,  13'd285,  -13'd404,  13'd332,  
-13'd252,  13'd520,  13'd434,  -13'd551,  -13'd736,  -13'd220,  13'd549,  -13'd93,  13'd1278,  13'd493,  -13'd83,  13'd341,  -13'd509,  13'd1,  13'd84,  -13'd598,  
-13'd8,  -13'd281,  -13'd9,  -13'd65,  -13'd179,  13'd238,  -13'd197,  -13'd493,  13'd569,  13'd677,  -13'd675,  -13'd419,  -13'd399,  13'd762,  -13'd316,  -13'd1193,  
-13'd146,  -13'd100,  -13'd654,  13'd120,  -13'd51,  -13'd317,  -13'd274,  -13'd49,  13'd494,  13'd309,  -13'd851,  13'd130,  -13'd369,  -13'd8,  -13'd414,  -13'd180,  
13'd228,  -13'd9,  -13'd239,  13'd240,  -13'd54,  13'd592,  -13'd852,  -13'd52,  13'd342,  -13'd106,  -13'd233,  -13'd643,  -13'd342,  -13'd313,  -13'd159,  -13'd626,  
13'd988,  -13'd281,  13'd360,  -13'd55,  -13'd1863,  13'd704,  -13'd480,  -13'd85,  13'd163,  -13'd357,  -13'd392,  13'd1214,  -13'd83,  13'd901,  13'd565,  -13'd355,  
13'd309,  -13'd193,  13'd525,  -13'd76,  -13'd67,  13'd448,  13'd1172,  13'd438,  -13'd48,  13'd431,  13'd172,  13'd190,  13'd145,  13'd620,  13'd581,  -13'd211,  
13'd14,  -13'd497,  -13'd263,  -13'd241,  13'd305,  -13'd336,  13'd176,  13'd410,  13'd415,  -13'd737,  13'd228,  -13'd699,  -13'd268,  13'd44,  -13'd123,  13'd82,  
-13'd21,  -13'd272,  13'd383,  13'd527,  -13'd306,  -13'd442,  13'd146,  13'd62,  -13'd196,  -13'd278,  13'd66,  -13'd733,  13'd326,  -13'd76,  -13'd574,  -13'd211,  
-13'd741,  -13'd700,  -13'd480,  -13'd58,  13'd224,  -13'd444,  13'd81,  -13'd152,  13'd199,  13'd848,  -13'd497,  -13'd112,  13'd639,  -13'd398,  -13'd543,  13'd429,  

13'd403,  13'd544,  -13'd588,  -13'd492,  13'd636,  -13'd516,  -13'd625,  13'd891,  -13'd329,  13'd296,  13'd11,  13'd87,  13'd618,  13'd67,  -13'd652,  13'd603,  
-13'd315,  -13'd363,  -13'd476,  13'd326,  13'd606,  -13'd361,  -13'd1025,  13'd667,  13'd115,  13'd73,  -13'd66,  13'd310,  13'd173,  13'd357,  13'd536,  13'd106,  
13'd589,  -13'd314,  -13'd153,  -13'd104,  -13'd620,  13'd565,  13'd321,  -13'd689,  13'd113,  -13'd635,  13'd1156,  13'd64,  13'd327,  13'd359,  -13'd72,  13'd567,  
-13'd435,  -13'd366,  -13'd325,  13'd169,  -13'd107,  13'd13,  13'd1023,  -13'd430,  -13'd431,  13'd119,  13'd203,  13'd182,  13'd505,  -13'd428,  13'd349,  -13'd236,  
-13'd178,  13'd79,  13'd32,  -13'd494,  -13'd566,  -13'd308,  13'd518,  13'd132,  -13'd340,  -13'd821,  13'd110,  -13'd456,  -13'd567,  13'd863,  13'd357,  13'd7,  
13'd15,  13'd78,  -13'd766,  -13'd58,  13'd116,  -13'd779,  -13'd877,  -13'd122,  -13'd310,  13'd264,  13'd833,  -13'd118,  -13'd146,  13'd86,  13'd74,  -13'd272,  
13'd630,  -13'd120,  13'd585,  13'd97,  13'd115,  -13'd442,  -13'd40,  -13'd711,  -13'd731,  13'd445,  13'd523,  13'd853,  13'd214,  -13'd220,  13'd308,  13'd344,  
-13'd272,  -13'd338,  13'd197,  13'd109,  13'd512,  -13'd959,  -13'd440,  13'd133,  -13'd499,  13'd967,  13'd951,  13'd544,  -13'd80,  -13'd3,  13'd438,  -13'd102,  
-13'd202,  -13'd38,  -13'd335,  -13'd585,  -13'd408,  -13'd1084,  13'd258,  -13'd245,  -13'd463,  13'd747,  13'd17,  -13'd264,  13'd720,  -13'd19,  -13'd355,  13'd196,  
-13'd458,  13'd652,  13'd596,  -13'd731,  13'd145,  -13'd55,  -13'd107,  13'd804,  -13'd860,  13'd1056,  -13'd322,  13'd527,  -13'd687,  13'd167,  -13'd869,  -13'd377,  
-13'd729,  -13'd676,  -13'd354,  -13'd644,  -13'd221,  13'd105,  -13'd506,  -13'd660,  13'd493,  13'd589,  13'd302,  -13'd84,  13'd148,  13'd289,  -13'd205,  13'd364,  
13'd98,  -13'd705,  -13'd188,  13'd531,  13'd124,  -13'd323,  -13'd1031,  -13'd136,  13'd236,  13'd330,  -13'd222,  13'd53,  -13'd372,  13'd163,  -13'd712,  13'd603,  
13'd345,  -13'd803,  13'd97,  13'd516,  13'd222,  -13'd29,  13'd43,  13'd113,  13'd727,  13'd927,  -13'd515,  13'd256,  -13'd404,  -13'd616,  -13'd499,  13'd317,  
-13'd1060,  13'd146,  -13'd196,  -13'd16,  13'd695,  -13'd158,  -13'd786,  13'd253,  13'd113,  13'd583,  -13'd475,  -13'd608,  13'd549,  -13'd202,  13'd613,  13'd625,  
-13'd331,  -13'd358,  -13'd744,  -13'd30,  13'd369,  13'd164,  -13'd103,  -13'd482,  13'd258,  13'd922,  -13'd73,  13'd649,  -13'd519,  13'd791,  13'd69,  -13'd639,  
-13'd395,  -13'd857,  13'd234,  -13'd203,  13'd344,  13'd38,  -13'd512,  -13'd422,  13'd904,  -13'd554,  13'd160,  -13'd556,  13'd468,  -13'd771,  13'd420,  13'd335,  
-13'd480,  -13'd577,  -13'd619,  -13'd148,  -13'd416,  13'd787,  -13'd779,  13'd411,  -13'd120,  13'd455,  13'd118,  13'd805,  13'd164,  -13'd510,  13'd173,  13'd107,  
13'd473,  -13'd315,  -13'd232,  13'd195,  -13'd398,  13'd700,  13'd225,  13'd637,  -13'd453,  -13'd527,  13'd667,  13'd496,  13'd10,  -13'd238,  -13'd13,  13'd35,  
-13'd7,  13'd801,  -13'd160,  13'd0,  13'd368,  -13'd30,  13'd115,  13'd650,  -13'd166,  13'd366,  -13'd116,  -13'd100,  -13'd201,  -13'd51,  -13'd89,  13'd113,  
-13'd41,  -13'd115,  13'd278,  -13'd27,  13'd824,  13'd107,  13'd103,  13'd875,  13'd581,  -13'd37,  13'd36,  -13'd750,  13'd154,  -13'd481,  13'd241,  13'd31,  
-13'd0,  -13'd285,  13'd400,  13'd552,  13'd181,  -13'd483,  13'd374,  -13'd187,  13'd310,  13'd195,  -13'd228,  13'd324,  13'd873,  13'd152,  13'd380,  13'd489,  
-13'd11,  -13'd204,  13'd24,  -13'd30,  -13'd655,  -13'd301,  13'd626,  13'd182,  13'd422,  -13'd926,  13'd288,  13'd216,  13'd531,  -13'd682,  13'd690,  13'd438,  
13'd728,  -13'd114,  -13'd587,  13'd271,  13'd307,  13'd191,  -13'd739,  -13'd42,  -13'd561,  13'd424,  13'd674,  13'd128,  13'd714,  -13'd461,  -13'd244,  -13'd431,  
13'd252,  13'd1087,  -13'd248,  13'd580,  -13'd24,  -13'd242,  -13'd286,  13'd208,  13'd72,  -13'd49,  -13'd95,  13'd701,  13'd245,  -13'd506,  13'd3,  -13'd300,  
13'd1013,  13'd727,  13'd399,  -13'd221,  -13'd65,  13'd286,  13'd178,  13'd93,  13'd997,  13'd1592,  -13'd560,  13'd1020,  13'd576,  13'd707,  13'd514,  13'd414,  

13'd668,  -13'd192,  -13'd857,  -13'd515,  13'd349,  -13'd62,  13'd357,  13'd272,  -13'd252,  13'd247,  13'd143,  -13'd314,  -13'd1092,  13'd265,  13'd464,  -13'd228,  
-13'd585,  13'd20,  -13'd1432,  13'd165,  13'd218,  13'd405,  13'd64,  -13'd76,  13'd446,  13'd106,  -13'd273,  13'd13,  -13'd748,  -13'd571,  -13'd353,  13'd222,  
-13'd58,  13'd154,  -13'd596,  13'd795,  -13'd289,  13'd821,  -13'd138,  -13'd80,  -13'd304,  13'd851,  13'd34,  13'd11,  13'd98,  -13'd956,  13'd492,  13'd88,  
-13'd464,  -13'd354,  -13'd324,  13'd418,  13'd107,  13'd62,  13'd49,  -13'd216,  13'd519,  13'd571,  -13'd226,  -13'd220,  13'd414,  -13'd508,  13'd107,  13'd606,  
-13'd346,  -13'd1084,  -13'd273,  13'd426,  13'd388,  13'd128,  -13'd93,  13'd154,  -13'd81,  13'd513,  13'd130,  -13'd243,  -13'd873,  13'd365,  -13'd11,  13'd260,  
13'd437,  13'd307,  -13'd302,  -13'd283,  13'd36,  13'd133,  -13'd217,  13'd438,  13'd447,  13'd7,  13'd29,  13'd89,  13'd74,  13'd37,  13'd110,  13'd485,  
13'd658,  13'd622,  -13'd52,  -13'd625,  -13'd338,  -13'd7,  -13'd680,  -13'd36,  13'd491,  13'd292,  -13'd1207,  -13'd337,  13'd156,  -13'd125,  13'd80,  13'd769,  
-13'd40,  -13'd172,  -13'd248,  -13'd293,  13'd299,  -13'd0,  13'd317,  -13'd234,  -13'd81,  13'd474,  13'd222,  13'd954,  -13'd138,  -13'd95,  13'd583,  13'd498,  
13'd262,  -13'd112,  -13'd1394,  13'd624,  -13'd48,  13'd471,  -13'd219,  -13'd426,  13'd388,  13'd61,  -13'd438,  -13'd221,  -13'd117,  -13'd276,  13'd460,  13'd589,  
-13'd873,  -13'd747,  -13'd613,  13'd790,  -13'd808,  13'd31,  -13'd134,  13'd107,  13'd86,  -13'd1179,  13'd283,  -13'd272,  13'd737,  13'd396,  -13'd195,  -13'd404,  
13'd87,  -13'd504,  13'd285,  13'd228,  13'd19,  -13'd422,  -13'd510,  13'd395,  13'd607,  13'd198,  -13'd1008,  13'd345,  13'd918,  -13'd153,  13'd565,  13'd334,  
-13'd74,  -13'd280,  13'd399,  -13'd327,  -13'd503,  -13'd205,  13'd12,  13'd204,  -13'd16,  -13'd101,  -13'd580,  13'd85,  13'd386,  13'd763,  13'd99,  -13'd432,  
13'd644,  13'd138,  -13'd626,  13'd765,  13'd97,  -13'd113,  -13'd352,  13'd150,  -13'd277,  -13'd306,  13'd787,  -13'd13,  -13'd214,  -13'd343,  13'd278,  13'd223,  
13'd332,  13'd95,  13'd278,  13'd202,  -13'd759,  13'd530,  -13'd95,  13'd430,  -13'd247,  -13'd842,  13'd628,  13'd250,  13'd708,  13'd82,  -13'd483,  13'd570,  
-13'd186,  13'd586,  -13'd143,  13'd63,  13'd3,  13'd875,  13'd732,  13'd0,  13'd501,  13'd472,  13'd439,  -13'd462,  13'd156,  13'd550,  -13'd707,  13'd324,  
-13'd37,  -13'd286,  -13'd475,  -13'd160,  13'd1007,  -13'd461,  -13'd701,  -13'd225,  -13'd235,  13'd519,  13'd662,  -13'd836,  -13'd30,  -13'd525,  13'd277,  -13'd365,  
-13'd514,  13'd566,  -13'd71,  -13'd104,  13'd211,  -13'd90,  -13'd888,  -13'd59,  -13'd138,  -13'd112,  -13'd529,  -13'd318,  -13'd74,  -13'd628,  -13'd504,  13'd502,  
13'd368,  -13'd378,  -13'd88,  -13'd176,  13'd121,  -13'd412,  13'd118,  -13'd2,  13'd435,  -13'd309,  13'd121,  13'd386,  -13'd916,  -13'd64,  -13'd33,  13'd448,  
13'd559,  13'd290,  -13'd362,  -13'd886,  -13'd354,  13'd107,  13'd333,  -13'd344,  -13'd204,  -13'd473,  13'd65,  13'd435,  -13'd455,  13'd266,  13'd105,  -13'd401,  
-13'd665,  13'd141,  -13'd513,  13'd437,  -13'd226,  -13'd443,  -13'd111,  13'd82,  -13'd406,  -13'd520,  13'd271,  -13'd340,  -13'd234,  13'd379,  13'd135,  -13'd543,  
-13'd158,  13'd264,  -13'd320,  -13'd260,  13'd768,  13'd729,  -13'd44,  -13'd240,  13'd896,  -13'd475,  13'd974,  13'd375,  13'd319,  -13'd646,  13'd656,  13'd481,  
-13'd246,  -13'd509,  -13'd481,  -13'd648,  13'd811,  -13'd656,  13'd114,  -13'd545,  -13'd106,  13'd284,  13'd105,  -13'd401,  -13'd227,  -13'd320,  -13'd171,  -13'd408,  
13'd174,  13'd462,  -13'd127,  -13'd309,  -13'd48,  -13'd197,  -13'd447,  -13'd1050,  13'd913,  13'd695,  -13'd115,  13'd562,  -13'd327,  13'd988,  13'd60,  -13'd210,  
-13'd133,  13'd211,  -13'd16,  -13'd187,  -13'd388,  -13'd284,  -13'd45,  -13'd562,  13'd88,  -13'd110,  -13'd33,  13'd89,  13'd61,  13'd954,  -13'd433,  13'd122,  
-13'd751,  -13'd110,  13'd681,  13'd381,  13'd8,  -13'd115,  13'd231,  13'd442,  13'd609,  -13'd418,  -13'd193,  -13'd754,  -13'd692,  -13'd73,  -13'd68,  -13'd720,  

13'd410,  13'd391,  13'd650,  -13'd662,  -13'd171,  13'd353,  13'd408,  13'd101,  13'd659,  13'd37,  -13'd689,  -13'd286,  13'd151,  -13'd82,  -13'd225,  13'd284,  
-13'd550,  13'd944,  13'd585,  13'd276,  13'd759,  13'd66,  -13'd316,  -13'd244,  -13'd766,  -13'd153,  -13'd1099,  13'd328,  13'd410,  -13'd284,  13'd366,  13'd346,  
13'd407,  -13'd319,  -13'd291,  13'd17,  -13'd388,  -13'd959,  13'd298,  -13'd250,  13'd228,  13'd107,  13'd12,  13'd314,  -13'd775,  13'd197,  13'd89,  13'd82,  
-13'd508,  -13'd655,  13'd780,  -13'd197,  -13'd228,  -13'd660,  -13'd153,  13'd164,  -13'd148,  -13'd576,  -13'd163,  -13'd460,  -13'd665,  13'd889,  13'd253,  13'd489,  
-13'd498,  13'd762,  13'd298,  13'd25,  -13'd378,  13'd199,  13'd192,  13'd55,  13'd747,  -13'd168,  -13'd99,  -13'd714,  -13'd537,  13'd822,  -13'd270,  13'd554,  
13'd127,  13'd387,  -13'd326,  -13'd386,  13'd360,  -13'd180,  13'd89,  13'd818,  -13'd362,  -13'd228,  -13'd647,  -13'd15,  -13'd838,  13'd171,  -13'd500,  13'd1,  
-13'd439,  -13'd300,  13'd98,  13'd103,  13'd687,  13'd235,  -13'd560,  13'd268,  -13'd172,  13'd424,  -13'd1130,  13'd299,  -13'd357,  -13'd948,  13'd271,  -13'd437,  
-13'd247,  -13'd394,  13'd89,  -13'd231,  13'd21,  13'd358,  -13'd165,  -13'd547,  13'd177,  13'd517,  13'd22,  -13'd158,  -13'd371,  -13'd370,  -13'd279,  -13'd489,  
-13'd488,  -13'd872,  13'd710,  -13'd80,  -13'd274,  -13'd557,  -13'd12,  13'd122,  -13'd395,  -13'd188,  13'd337,  13'd90,  -13'd540,  13'd562,  13'd495,  -13'd458,  
-13'd516,  13'd108,  -13'd253,  -13'd215,  -13'd54,  13'd259,  -13'd63,  13'd998,  -13'd33,  13'd225,  -13'd214,  13'd160,  13'd316,  13'd438,  -13'd616,  -13'd1075,  
13'd20,  -13'd140,  13'd161,  -13'd320,  13'd794,  -13'd1,  -13'd560,  13'd3,  13'd485,  13'd19,  -13'd720,  13'd190,  13'd537,  -13'd593,  -13'd479,  13'd20,  
13'd223,  13'd727,  13'd499,  13'd380,  -13'd500,  13'd435,  -13'd418,  13'd262,  -13'd406,  13'd666,  13'd757,  13'd356,  13'd480,  -13'd682,  13'd139,  13'd774,  
-13'd46,  -13'd531,  -13'd9,  13'd662,  13'd227,  13'd759,  -13'd338,  13'd963,  -13'd468,  -13'd376,  13'd925,  13'd448,  13'd613,  -13'd343,  -13'd301,  -13'd59,  
13'd63,  -13'd272,  -13'd222,  -13'd387,  -13'd453,  -13'd553,  13'd541,  -13'd705,  13'd706,  -13'd150,  13'd805,  -13'd37,  13'd221,  -13'd9,  -13'd387,  -13'd290,  
13'd332,  -13'd315,  -13'd1081,  13'd544,  -13'd200,  13'd445,  13'd24,  13'd414,  13'd233,  -13'd358,  -13'd113,  13'd130,  13'd593,  -13'd507,  13'd382,  13'd531,  
13'd98,  -13'd714,  -13'd635,  13'd187,  13'd202,  13'd83,  13'd572,  13'd361,  13'd8,  13'd110,  13'd1272,  13'd102,  13'd785,  13'd766,  13'd602,  13'd260,  
13'd509,  -13'd753,  13'd665,  13'd236,  13'd170,  13'd557,  13'd274,  -13'd127,  -13'd480,  13'd230,  -13'd81,  -13'd84,  13'd678,  13'd113,  13'd324,  13'd384,  
13'd15,  13'd731,  13'd731,  13'd544,  13'd150,  13'd255,  -13'd23,  -13'd418,  -13'd206,  -13'd147,  13'd690,  13'd31,  -13'd490,  -13'd422,  -13'd368,  13'd495,  
13'd63,  13'd366,  13'd145,  13'd121,  13'd937,  13'd100,  -13'd164,  -13'd30,  -13'd238,  -13'd232,  13'd291,  13'd61,  13'd145,  13'd92,  -13'd373,  -13'd446,  
13'd693,  -13'd146,  -13'd197,  13'd762,  -13'd707,  13'd423,  13'd80,  -13'd76,  13'd250,  13'd481,  -13'd42,  13'd164,  -13'd118,  13'd244,  -13'd66,  -13'd509,  
13'd439,  13'd505,  13'd553,  13'd153,  -13'd652,  -13'd67,  -13'd27,  -13'd12,  -13'd440,  13'd349,  13'd661,  -13'd560,  13'd696,  13'd475,  13'd217,  -13'd72,  
-13'd172,  13'd203,  -13'd434,  -13'd153,  -13'd83,  -13'd220,  13'd519,  -13'd146,  -13'd320,  -13'd94,  -13'd300,  -13'd55,  13'd755,  13'd284,  -13'd47,  -13'd181,  
13'd490,  13'd369,  13'd329,  13'd451,  -13'd3,  13'd364,  -13'd320,  -13'd390,  13'd516,  -13'd346,  13'd296,  -13'd271,  -13'd170,  -13'd189,  -13'd258,  -13'd74,  
-13'd697,  13'd797,  13'd457,  -13'd89,  -13'd430,  -13'd196,  -13'd346,  13'd473,  13'd450,  -13'd30,  -13'd358,  -13'd11,  -13'd147,  13'd480,  13'd475,  13'd847,  
13'd890,  13'd101,  13'd847,  13'd368,  13'd202,  -13'd124,  13'd418,  13'd530,  13'd635,  13'd133,  13'd268,  13'd773,  -13'd325,  13'd92,  13'd846,  13'd405,  

13'd38,  13'd207,  13'd950,  -13'd272,  -13'd931,  -13'd172,  13'd854,  -13'd427,  -13'd264,  -13'd807,  13'd231,  -13'd253,  -13'd573,  13'd894,  13'd414,  13'd56,  
-13'd358,  -13'd223,  13'd324,  -13'd5,  13'd515,  -13'd237,  13'd1065,  -13'd1016,  13'd378,  -13'd366,  13'd1448,  -13'd290,  -13'd401,  13'd203,  -13'd526,  -13'd484,  
13'd180,  13'd78,  13'd54,  -13'd843,  -13'd21,  -13'd781,  -13'd64,  -13'd869,  13'd490,  13'd353,  13'd436,  13'd239,  13'd352,  13'd1214,  -13'd350,  -13'd569,  
13'd481,  13'd451,  -13'd687,  -13'd145,  -13'd598,  -13'd274,  13'd371,  13'd319,  13'd611,  -13'd283,  13'd219,  -13'd653,  -13'd155,  -13'd675,  -13'd85,  -13'd326,  
13'd971,  13'd409,  -13'd389,  13'd919,  -13'd221,  13'd120,  -13'd481,  13'd348,  -13'd81,  -13'd154,  -13'd86,  13'd645,  13'd878,  13'd999,  13'd253,  13'd887,  
-13'd23,  13'd350,  13'd231,  -13'd452,  13'd10,  13'd221,  13'd814,  -13'd23,  -13'd740,  -13'd386,  -13'd383,  13'd609,  -13'd459,  13'd469,  -13'd193,  -13'd497,  
13'd393,  -13'd732,  -13'd178,  -13'd120,  -13'd85,  -13'd327,  13'd613,  13'd289,  13'd451,  -13'd652,  -13'd186,  13'd588,  13'd56,  13'd108,  13'd37,  -13'd259,  
-13'd64,  -13'd276,  13'd92,  13'd561,  13'd256,  -13'd75,  -13'd552,  -13'd902,  13'd623,  13'd1191,  13'd656,  -13'd28,  -13'd466,  13'd289,  -13'd271,  -13'd406,  
-13'd85,  -13'd392,  -13'd1538,  -13'd677,  -13'd49,  -13'd289,  -13'd824,  13'd360,  -13'd55,  13'd489,  13'd158,  -13'd938,  13'd646,  -13'd737,  -13'd467,  13'd256,  
-13'd777,  -13'd39,  -13'd403,  13'd194,  13'd543,  13'd624,  -13'd661,  -13'd155,  -13'd605,  13'd997,  13'd399,  13'd108,  13'd603,  -13'd506,  -13'd151,  13'd287,  
13'd75,  -13'd115,  13'd461,  13'd507,  -13'd312,  -13'd102,  13'd270,  -13'd250,  13'd489,  13'd184,  -13'd181,  13'd124,  13'd395,  13'd512,  13'd839,  13'd464,  
13'd208,  -13'd427,  13'd702,  13'd913,  -13'd273,  13'd223,  -13'd430,  13'd976,  -13'd103,  13'd177,  13'd46,  -13'd425,  13'd880,  13'd787,  13'd573,  -13'd550,  
-13'd207,  -13'd612,  -13'd228,  13'd352,  13'd810,  13'd75,  13'd251,  -13'd704,  -13'd35,  13'd91,  13'd540,  13'd254,  13'd177,  -13'd719,  13'd27,  -13'd482,  
-13'd332,  -13'd292,  -13'd1299,  -13'd181,  -13'd34,  13'd286,  -13'd377,  -13'd199,  13'd519,  -13'd630,  13'd382,  13'd43,  13'd174,  -13'd698,  -13'd476,  -13'd251,  
-13'd864,  13'd7,  -13'd282,  13'd1047,  -13'd97,  13'd246,  -13'd930,  13'd393,  13'd114,  13'd530,  13'd889,  -13'd344,  13'd286,  -13'd82,  13'd216,  -13'd285,  
13'd111,  13'd71,  13'd356,  13'd5,  -13'd18,  13'd445,  13'd176,  -13'd319,  -13'd489,  -13'd21,  -13'd66,  13'd135,  13'd385,  13'd157,  -13'd177,  -13'd122,  
13'd17,  -13'd338,  13'd79,  13'd516,  13'd510,  -13'd647,  -13'd1200,  -13'd189,  -13'd641,  -13'd101,  -13'd289,  13'd191,  13'd166,  13'd173,  13'd197,  13'd301,  
13'd657,  13'd122,  13'd933,  -13'd80,  13'd354,  13'd20,  13'd633,  -13'd279,  -13'd396,  13'd95,  -13'd108,  13'd836,  13'd628,  13'd477,  13'd2,  13'd145,  
13'd129,  -13'd39,  13'd36,  -13'd220,  13'd1121,  13'd48,  13'd100,  -13'd172,  13'd332,  -13'd482,  13'd820,  13'd523,  -13'd226,  13'd253,  -13'd57,  -13'd220,  
-13'd3,  13'd379,  13'd199,  -13'd92,  13'd352,  13'd97,  13'd23,  13'd484,  13'd138,  -13'd204,  -13'd374,  -13'd461,  -13'd857,  13'd414,  -13'd63,  -13'd557,  
13'd584,  13'd99,  -13'd240,  -13'd301,  -13'd125,  13'd65,  13'd665,  13'd62,  13'd552,  13'd144,  -13'd90,  13'd50,  13'd241,  -13'd139,  -13'd400,  13'd277,  
-13'd366,  -13'd313,  13'd39,  -13'd100,  -13'd357,  -13'd210,  -13'd383,  -13'd459,  13'd479,  13'd251,  13'd710,  -13'd86,  13'd397,  -13'd1173,  13'd394,  13'd358,  
-13'd385,  13'd180,  13'd522,  13'd96,  -13'd400,  -13'd805,  13'd270,  -13'd129,  13'd441,  13'd464,  13'd191,  13'd126,  -13'd175,  13'd677,  13'd25,  13'd170,  
-13'd528,  13'd117,  13'd619,  -13'd338,  -13'd500,  -13'd200,  -13'd134,  13'd470,  13'd279,  -13'd359,  -13'd704,  -13'd86,  13'd428,  13'd123,  13'd248,  -13'd227,  
-13'd364,  13'd187,  13'd6,  -13'd58,  -13'd677,  13'd199,  -13'd330,  13'd471,  -13'd325,  -13'd754,  -13'd369,  -13'd624,  -13'd25,  13'd740,  13'd386,  -13'd662,  

-13'd1,  13'd339,  -13'd240,  13'd125,  -13'd761,  -13'd274,  13'd512,  13'd314,  13'd391,  13'd17,  -13'd264,  -13'd50,  -13'd254,  -13'd332,  13'd862,  13'd147,  
-13'd81,  13'd315,  -13'd47,  13'd306,  -13'd38,  13'd441,  -13'd349,  13'd490,  13'd409,  13'd409,  13'd892,  -13'd453,  -13'd681,  -13'd948,  13'd231,  13'd193,  
13'd350,  13'd305,  -13'd358,  13'd259,  13'd174,  13'd262,  -13'd1092,  -13'd0,  13'd114,  13'd25,  13'd687,  -13'd64,  13'd517,  -13'd1318,  13'd160,  -13'd171,  
13'd33,  -13'd283,  13'd356,  -13'd30,  -13'd421,  13'd365,  -13'd863,  13'd344,  -13'd86,  13'd144,  -13'd325,  -13'd55,  13'd87,  -13'd1895,  -13'd69,  13'd286,  
-13'd688,  -13'd788,  13'd159,  -13'd429,  -13'd200,  -13'd422,  -13'd490,  -13'd51,  13'd276,  13'd267,  -13'd162,  13'd372,  -13'd327,  13'd150,  -13'd327,  13'd15,  
-13'd34,  -13'd487,  13'd1048,  13'd852,  -13'd184,  13'd250,  -13'd388,  13'd351,  -13'd104,  -13'd33,  13'd131,  13'd341,  13'd402,  -13'd350,  13'd18,  13'd221,  
-13'd769,  -13'd358,  -13'd149,  -13'd66,  13'd301,  13'd557,  13'd574,  13'd241,  13'd229,  -13'd97,  -13'd145,  13'd104,  -13'd401,  -13'd423,  -13'd58,  13'd168,  
-13'd1084,  -13'd128,  -13'd758,  13'd719,  13'd350,  13'd504,  -13'd854,  -13'd241,  -13'd372,  -13'd106,  -13'd247,  -13'd450,  -13'd470,  -13'd736,  -13'd160,  -13'd463,  
-13'd581,  13'd468,  13'd1,  -13'd605,  13'd508,  13'd42,  -13'd434,  -13'd604,  -13'd722,  13'd760,  -13'd430,  -13'd664,  -13'd222,  -13'd321,  13'd99,  13'd308,  
-13'd1275,  -13'd109,  13'd136,  -13'd88,  -13'd355,  -13'd357,  13'd268,  13'd67,  13'd205,  13'd380,  13'd169,  -13'd908,  -13'd271,  13'd78,  -13'd139,  -13'd613,  
13'd92,  13'd167,  13'd352,  13'd517,  13'd421,  13'd215,  -13'd69,  13'd465,  -13'd936,  13'd5,  13'd324,  13'd482,  13'd528,  13'd451,  13'd211,  13'd177,  
-13'd737,  13'd327,  -13'd399,  13'd115,  13'd870,  -13'd105,  -13'd247,  13'd84,  13'd946,  13'd158,  13'd493,  13'd447,  13'd99,  -13'd987,  -13'd117,  -13'd197,  
13'd143,  13'd300,  13'd56,  -13'd219,  13'd855,  13'd58,  13'd19,  13'd183,  13'd11,  13'd238,  13'd188,  13'd416,  -13'd613,  13'd386,  -13'd352,  13'd617,  
13'd373,  -13'd701,  13'd699,  -13'd117,  -13'd591,  -13'd133,  -13'd152,  -13'd42,  -13'd434,  -13'd924,  13'd370,  -13'd49,  13'd120,  13'd424,  13'd501,  -13'd162,  
13'd563,  -13'd595,  13'd704,  -13'd522,  -13'd134,  13'd826,  -13'd154,  13'd154,  13'd530,  13'd161,  -13'd83,  -13'd121,  13'd63,  13'd459,  -13'd13,  13'd328,  
13'd1023,  13'd25,  13'd102,  -13'd581,  -13'd527,  -13'd282,  13'd435,  -13'd437,  13'd601,  -13'd46,  13'd499,  13'd757,  -13'd572,  -13'd615,  13'd15,  -13'd458,  
-13'd39,  -13'd165,  -13'd771,  13'd208,  -13'd99,  -13'd185,  -13'd80,  -13'd540,  13'd905,  -13'd270,  13'd44,  13'd746,  13'd447,  13'd330,  -13'd615,  13'd598,  
13'd373,  -13'd337,  -13'd172,  13'd14,  -13'd440,  13'd552,  13'd543,  -13'd293,  13'd301,  -13'd194,  -13'd533,  13'd167,  13'd430,  -13'd275,  -13'd378,  13'd244,  
13'd583,  13'd345,  13'd767,  13'd393,  13'd534,  -13'd358,  13'd74,  13'd233,  -13'd45,  -13'd215,  13'd250,  -13'd786,  13'd397,  13'd1,  13'd398,  13'd27,  
-13'd583,  13'd657,  -13'd474,  -13'd142,  -13'd121,  -13'd632,  -13'd437,  -13'd133,  -13'd255,  13'd952,  13'd150,  13'd110,  13'd742,  -13'd83,  13'd227,  -13'd416,  
13'd718,  13'd609,  13'd170,  -13'd178,  13'd217,  -13'd23,  13'd1277,  -13'd186,  -13'd237,  -13'd788,  13'd163,  13'd609,  -13'd502,  -13'd248,  -13'd708,  13'd300,  
13'd56,  13'd203,  -13'd703,  -13'd267,  -13'd244,  -13'd134,  13'd1415,  -13'd284,  13'd773,  13'd291,  13'd301,  -13'd198,  -13'd302,  13'd567,  -13'd727,  -13'd625,  
13'd119,  -13'd273,  13'd453,  -13'd147,  13'd16,  -13'd324,  -13'd102,  -13'd162,  13'd281,  13'd54,  -13'd62,  -13'd720,  13'd456,  13'd681,  -13'd285,  -13'd560,  
-13'd60,  13'd753,  13'd90,  -13'd246,  -13'd195,  13'd910,  -13'd167,  13'd221,  -13'd61,  13'd407,  13'd159,  -13'd345,  13'd236,  -13'd398,  13'd37,  13'd193,  
-13'd1092,  -13'd930,  -13'd876,  13'd642,  13'd123,  13'd565,  13'd269,  -13'd280,  -13'd405,  13'd680,  -13'd477,  -13'd766,  -13'd343,  -13'd775,  13'd544,  -13'd236,  

13'd587,  13'd187,  13'd52,  13'd96,  -13'd312,  13'd187,  13'd881,  13'd214,  13'd218,  -13'd208,  13'd438,  13'd304,  13'd45,  13'd369,  -13'd60,  13'd238,  
13'd256,  13'd369,  13'd638,  13'd323,  13'd347,  13'd210,  13'd122,  -13'd33,  13'd463,  13'd425,  13'd1028,  13'd126,  13'd145,  13'd538,  -13'd23,  -13'd368,  
-13'd359,  -13'd814,  13'd346,  -13'd98,  13'd99,  13'd468,  13'd703,  13'd745,  -13'd135,  13'd499,  13'd425,  13'd352,  13'd171,  -13'd331,  13'd433,  13'd321,  
-13'd109,  -13'd422,  13'd371,  13'd295,  -13'd562,  -13'd96,  -13'd113,  -13'd102,  -13'd249,  13'd611,  -13'd622,  -13'd37,  13'd551,  -13'd184,  -13'd370,  13'd5,  
-13'd309,  -13'd270,  -13'd643,  -13'd559,  -13'd25,  -13'd391,  -13'd79,  -13'd34,  -13'd317,  13'd82,  13'd16,  -13'd355,  13'd354,  13'd117,  -13'd239,  -13'd265,  
-13'd20,  13'd492,  -13'd211,  13'd372,  13'd221,  13'd578,  -13'd254,  -13'd64,  13'd270,  13'd441,  -13'd64,  -13'd378,  -13'd503,  13'd650,  13'd74,  -13'd555,  
-13'd188,  13'd45,  13'd562,  -13'd508,  -13'd324,  -13'd627,  -13'd44,  13'd90,  13'd225,  13'd79,  13'd514,  13'd56,  -13'd69,  13'd653,  13'd99,  13'd487,  
-13'd73,  -13'd698,  13'd28,  13'd277,  -13'd120,  13'd421,  -13'd55,  13'd222,  13'd9,  13'd188,  -13'd597,  -13'd264,  13'd535,  13'd421,  13'd167,  13'd216,  
-13'd243,  -13'd899,  13'd3,  13'd351,  13'd402,  13'd273,  -13'd97,  13'd240,  -13'd132,  -13'd368,  -13'd268,  -13'd597,  -13'd128,  13'd51,  -13'd105,  13'd23,  
-13'd1617,  -13'd588,  -13'd808,  -13'd325,  -13'd548,  -13'd1183,  -13'd59,  -13'd162,  -13'd995,  -13'd104,  -13'd52,  13'd288,  -13'd872,  13'd317,  -13'd468,  -13'd264,  
-13'd715,  -13'd784,  13'd743,  -13'd154,  13'd273,  13'd290,  -13'd380,  13'd586,  13'd342,  13'd688,  -13'd733,  -13'd133,  13'd49,  13'd1145,  13'd510,  -13'd103,  
13'd31,  -13'd221,  13'd353,  13'd488,  -13'd102,  -13'd192,  -13'd673,  -13'd94,  -13'd706,  -13'd830,  -13'd69,  13'd9,  13'd229,  13'd31,  13'd787,  13'd191,  
13'd46,  -13'd196,  13'd483,  13'd403,  -13'd607,  13'd258,  -13'd977,  -13'd363,  13'd376,  13'd301,  -13'd222,  -13'd480,  13'd55,  -13'd476,  13'd102,  -13'd66,  
13'd193,  -13'd416,  -13'd167,  -13'd345,  -13'd117,  13'd333,  -13'd387,  -13'd451,  -13'd508,  -13'd308,  -13'd579,  -13'd270,  -13'd494,  13'd236,  13'd98,  -13'd741,  
-13'd7,  -13'd288,  13'd70,  13'd67,  -13'd635,  13'd151,  13'd130,  13'd149,  13'd151,  13'd609,  -13'd281,  13'd103,  -13'd821,  -13'd292,  -13'd632,  13'd197,  
-13'd816,  13'd231,  -13'd294,  -13'd108,  13'd705,  13'd231,  -13'd693,  13'd679,  13'd56,  13'd693,  -13'd740,  -13'd66,  13'd74,  13'd121,  -13'd597,  -13'd432,  
-13'd482,  13'd678,  13'd326,  -13'd135,  -13'd591,  13'd52,  -13'd1068,  13'd29,  13'd264,  -13'd242,  13'd511,  13'd123,  -13'd551,  -13'd401,  -13'd150,  -13'd188,  
-13'd659,  -13'd168,  13'd75,  -13'd647,  13'd32,  -13'd846,  13'd418,  13'd216,  -13'd865,  -13'd159,  -13'd291,  13'd469,  13'd237,  13'd63,  -13'd181,  13'd692,  
13'd174,  13'd178,  13'd39,  13'd121,  -13'd590,  -13'd288,  13'd37,  13'd22,  13'd607,  13'd89,  -13'd224,  13'd825,  13'd57,  13'd509,  13'd767,  -13'd172,  
-13'd443,  13'd214,  13'd352,  -13'd785,  -13'd684,  13'd291,  13'd704,  13'd292,  -13'd560,  13'd647,  13'd6,  13'd14,  -13'd321,  -13'd361,  13'd432,  -13'd812,  
-13'd999,  13'd188,  -13'd827,  13'd252,  13'd844,  -13'd612,  13'd447,  -13'd290,  13'd1071,  -13'd151,  -13'd17,  -13'd331,  -13'd326,  -13'd312,  -13'd183,  -13'd232,  
-13'd22,  -13'd224,  -13'd680,  -13'd154,  13'd896,  13'd439,  13'd173,  -13'd937,  13'd330,  13'd247,  13'd559,  13'd55,  -13'd312,  -13'd813,  -13'd19,  13'd541,  
13'd512,  13'd557,  -13'd165,  13'd0,  -13'd274,  -13'd344,  -13'd173,  -13'd317,  13'd501,  13'd161,  13'd248,  13'd436,  13'd211,  13'd332,  -13'd157,  -13'd474,  
13'd612,  13'd344,  13'd428,  13'd247,  13'd591,  13'd1026,  13'd367,  13'd487,  -13'd229,  13'd173,  -13'd86,  13'd495,  13'd829,  -13'd6,  13'd11,  13'd387,  
13'd425,  -13'd288,  13'd757,  -13'd12,  13'd166,  13'd315,  13'd623,  13'd486,  13'd155,  -13'd599,  -13'd7,  13'd750,  13'd166,  13'd5,  13'd62,  -13'd173,  

13'd860,  13'd79,  13'd906,  13'd269,  13'd14,  13'd447,  13'd175,  -13'd842,  -13'd177,  13'd271,  13'd305,  13'd303,  -13'd143,  -13'd380,  13'd138,  -13'd74,  
-13'd44,  13'd408,  13'd778,  -13'd14,  -13'd12,  13'd365,  -13'd138,  -13'd229,  13'd40,  -13'd389,  -13'd390,  13'd197,  -13'd183,  -13'd133,  -13'd5,  13'd297,  
13'd101,  13'd86,  -13'd649,  13'd273,  13'd155,  13'd63,  13'd139,  13'd433,  13'd510,  -13'd227,  13'd137,  13'd38,  -13'd649,  13'd186,  -13'd356,  13'd297,  
13'd82,  -13'd310,  13'd294,  -13'd948,  13'd135,  -13'd83,  13'd185,  -13'd240,  13'd677,  13'd69,  13'd138,  13'd698,  -13'd655,  13'd1510,  -13'd522,  -13'd527,  
-13'd206,  13'd160,  13'd549,  13'd346,  13'd17,  13'd142,  13'd153,  -13'd29,  13'd416,  -13'd63,  -13'd47,  -13'd138,  -13'd414,  13'd966,  -13'd473,  -13'd268,  
-13'd123,  13'd631,  -13'd367,  -13'd301,  -13'd261,  13'd665,  13'd308,  -13'd138,  -13'd108,  13'd15,  13'd79,  -13'd115,  -13'd308,  13'd129,  13'd160,  13'd55,  
-13'd22,  -13'd161,  13'd683,  -13'd630,  -13'd108,  13'd573,  13'd147,  13'd422,  -13'd290,  13'd21,  -13'd479,  -13'd25,  -13'd269,  13'd447,  13'd955,  -13'd267,  
13'd1210,  -13'd584,  13'd830,  13'd381,  13'd378,  13'd18,  13'd733,  -13'd121,  -13'd100,  13'd71,  -13'd202,  13'd564,  -13'd220,  -13'd4,  13'd183,  -13'd822,  
-13'd78,  -13'd616,  -13'd69,  13'd474,  13'd307,  13'd37,  13'd276,  -13'd669,  13'd129,  -13'd209,  -13'd822,  13'd19,  13'd610,  13'd772,  -13'd395,  -13'd207,  
13'd183,  -13'd57,  -13'd361,  13'd355,  13'd913,  13'd628,  13'd538,  13'd175,  13'd381,  -13'd329,  -13'd439,  -13'd482,  13'd102,  13'd764,  -13'd1019,  -13'd334,  
-13'd165,  13'd758,  13'd5,  13'd112,  13'd56,  -13'd189,  13'd686,  13'd164,  -13'd352,  -13'd267,  13'd32,  -13'd517,  13'd226,  -13'd175,  -13'd380,  13'd506,  
-13'd210,  -13'd361,  13'd327,  13'd478,  13'd768,  13'd734,  13'd557,  13'd357,  13'd240,  -13'd550,  -13'd670,  -13'd602,  13'd428,  13'd508,  -13'd466,  13'd24,  
13'd667,  13'd408,  -13'd216,  -13'd51,  -13'd34,  13'd847,  -13'd386,  13'd192,  13'd424,  -13'd666,  -13'd375,  13'd192,  13'd349,  -13'd804,  13'd837,  -13'd670,  
13'd65,  -13'd79,  13'd138,  -13'd244,  -13'd7,  13'd89,  13'd152,  -13'd458,  -13'd315,  13'd161,  -13'd149,  13'd66,  -13'd33,  13'd212,  13'd518,  13'd347,  
13'd321,  -13'd951,  -13'd355,  -13'd179,  13'd733,  13'd294,  13'd693,  13'd214,  -13'd304,  13'd294,  -13'd589,  -13'd509,  -13'd83,  13'd953,  13'd98,  13'd184,  
13'd574,  13'd375,  13'd340,  13'd402,  -13'd653,  -13'd222,  13'd416,  13'd290,  13'd132,  -13'd19,  -13'd28,  -13'd28,  -13'd89,  13'd396,  -13'd288,  13'd320,  
13'd584,  -13'd140,  13'd97,  13'd261,  13'd1253,  -13'd177,  13'd358,  13'd264,  13'd629,  13'd23,  -13'd376,  -13'd310,  -13'd21,  13'd905,  -13'd191,  13'd113,  
13'd110,  13'd209,  -13'd103,  13'd32,  13'd350,  13'd32,  -13'd323,  -13'd458,  -13'd239,  -13'd432,  -13'd744,  13'd113,  -13'd661,  13'd682,  -13'd43,  13'd354,  
-13'd1,  -13'd799,  13'd411,  -13'd352,  -13'd273,  13'd114,  13'd21,  13'd134,  13'd530,  -13'd670,  -13'd459,  13'd314,  -13'd315,  -13'd123,  13'd300,  13'd192,  
-13'd652,  13'd52,  -13'd33,  13'd49,  -13'd440,  13'd8,  13'd933,  13'd11,  13'd612,  -13'd764,  -13'd78,  -13'd273,  -13'd61,  -13'd611,  -13'd5,  13'd175,  
13'd255,  13'd63,  -13'd136,  13'd350,  -13'd18,  -13'd689,  -13'd743,  -13'd120,  -13'd629,  13'd297,  -13'd1019,  -13'd644,  13'd4,  13'd589,  -13'd60,  13'd183,  
-13'd269,  13'd770,  13'd131,  13'd281,  13'd362,  -13'd201,  -13'd426,  13'd110,  -13'd554,  13'd23,  -13'd778,  -13'd383,  -13'd129,  13'd671,  13'd598,  13'd112,  
13'd466,  13'd539,  13'd185,  -13'd576,  -13'd90,  13'd100,  13'd35,  13'd461,  -13'd13,  -13'd492,  -13'd522,  -13'd520,  -13'd462,  13'd874,  13'd1194,  -13'd345,  
13'd265,  -13'd424,  13'd229,  13'd46,  13'd568,  -13'd377,  13'd597,  13'd604,  -13'd273,  -13'd934,  -13'd341,  -13'd497,  13'd295,  13'd1109,  13'd380,  13'd702,  
13'd86,  13'd570,  -13'd60,  13'd412,  13'd1058,  13'd728,  13'd271,  13'd336,  -13'd317,  -13'd913,  13'd94,  -13'd165,  -13'd379,  13'd512,  13'd56,  -13'd531,  

13'd485,  -13'd504,  -13'd867,  13'd29,  -13'd202,  13'd32,  -13'd581,  -13'd34,  -13'd43,  13'd482,  -13'd893,  -13'd29,  13'd652,  13'd117,  13'd840,  13'd278,  
-13'd87,  13'd232,  13'd343,  13'd219,  -13'd188,  13'd24,  -13'd1018,  13'd1038,  13'd445,  13'd701,  13'd105,  -13'd120,  -13'd169,  -13'd78,  13'd481,  13'd254,  
-13'd7,  -13'd707,  13'd502,  13'd155,  -13'd477,  13'd69,  -13'd93,  13'd528,  13'd218,  13'd58,  13'd1,  13'd544,  -13'd193,  -13'd240,  13'd553,  13'd118,  
13'd180,  13'd168,  13'd826,  13'd192,  -13'd807,  -13'd581,  -13'd882,  13'd36,  13'd75,  13'd438,  -13'd356,  13'd322,  13'd587,  -13'd838,  13'd470,  -13'd537,  
13'd361,  13'd592,  13'd121,  13'd513,  -13'd414,  -13'd193,  13'd111,  13'd600,  13'd96,  13'd394,  -13'd22,  13'd107,  13'd519,  -13'd634,  13'd165,  13'd574,  
13'd48,  13'd560,  -13'd117,  13'd807,  13'd109,  13'd486,  -13'd1009,  -13'd537,  13'd571,  13'd841,  -13'd648,  13'd109,  13'd500,  -13'd357,  13'd344,  -13'd548,  
-13'd468,  13'd76,  13'd311,  13'd685,  -13'd287,  13'd56,  -13'd180,  13'd0,  13'd238,  13'd799,  -13'd384,  -13'd490,  13'd428,  13'd823,  13'd331,  13'd147,  
13'd17,  13'd491,  13'd893,  13'd363,  13'd170,  -13'd704,  13'd54,  -13'd384,  13'd301,  -13'd56,  13'd584,  -13'd116,  13'd467,  13'd963,  -13'd306,  13'd745,  
-13'd484,  13'd691,  13'd337,  -13'd218,  -13'd291,  13'd453,  -13'd118,  13'd262,  -13'd507,  -13'd216,  13'd412,  13'd338,  -13'd106,  13'd179,  13'd140,  -13'd388,  
13'd677,  -13'd361,  13'd290,  13'd118,  -13'd631,  13'd477,  13'd240,  13'd322,  -13'd202,  -13'd325,  13'd106,  13'd851,  13'd202,  -13'd640,  -13'd283,  -13'd564,  
-13'd465,  13'd511,  -13'd33,  13'd62,  13'd600,  -13'd100,  -13'd927,  13'd745,  -13'd768,  -13'd176,  -13'd195,  13'd114,  -13'd431,  13'd177,  13'd36,  -13'd12,  
13'd49,  13'd315,  13'd154,  -13'd202,  13'd747,  13'd33,  13'd717,  -13'd106,  13'd134,  13'd283,  13'd175,  13'd117,  13'd14,  -13'd559,  -13'd251,  13'd105,  
-13'd478,  -13'd726,  13'd666,  -13'd566,  13'd468,  13'd442,  13'd286,  13'd160,  13'd113,  13'd178,  13'd322,  13'd340,  -13'd840,  13'd999,  13'd36,  -13'd614,  
13'd224,  -13'd382,  -13'd304,  13'd725,  13'd338,  -13'd816,  -13'd97,  13'd669,  13'd177,  13'd40,  -13'd257,  -13'd337,  -13'd0,  -13'd144,  13'd224,  -13'd54,  
13'd934,  13'd772,  13'd11,  -13'd463,  13'd28,  -13'd579,  -13'd101,  13'd289,  -13'd92,  -13'd815,  -13'd505,  -13'd193,  -13'd91,  13'd84,  13'd727,  13'd421,  
13'd340,  -13'd354,  -13'd193,  -13'd287,  -13'd177,  -13'd954,  13'd303,  -13'd645,  13'd248,  -13'd225,  -13'd478,  13'd930,  13'd193,  -13'd415,  -13'd380,  -13'd38,  
13'd795,  13'd357,  13'd136,  -13'd35,  -13'd148,  13'd136,  13'd1810,  -13'd301,  13'd1240,  -13'd49,  13'd291,  13'd36,  13'd416,  13'd948,  -13'd63,  13'd270,  
-13'd428,  13'd180,  -13'd116,  13'd127,  13'd151,  13'd552,  -13'd89,  -13'd388,  13'd476,  -13'd525,  13'd250,  -13'd304,  -13'd20,  13'd67,  -13'd353,  13'd209,  
-13'd731,  -13'd91,  -13'd418,  13'd213,  -13'd111,  -13'd559,  13'd324,  -13'd925,  13'd160,  13'd794,  -13'd387,  -13'd906,  -13'd512,  -13'd473,  -13'd70,  -13'd671,  
-13'd394,  13'd25,  -13'd99,  -13'd90,  13'd151,  -13'd288,  13'd85,  -13'd119,  -13'd263,  13'd713,  -13'd68,  13'd96,  -13'd411,  -13'd731,  13'd74,  13'd613,  
13'd198,  -13'd172,  13'd906,  -13'd245,  -13'd309,  -13'd215,  13'd731,  13'd28,  13'd168,  13'd285,  -13'd7,  -13'd380,  13'd499,  13'd1012,  -13'd366,  13'd280,  
-13'd87,  13'd103,  13'd338,  13'd318,  -13'd207,  13'd187,  -13'd429,  13'd424,  -13'd979,  -13'd373,  -13'd271,  -13'd71,  -13'd25,  13'd843,  -13'd53,  13'd100,  
13'd623,  -13'd598,  -13'd454,  -13'd599,  -13'd652,  -13'd560,  -13'd790,  13'd112,  -13'd905,  -13'd675,  13'd410,  -13'd179,  -13'd158,  -13'd25,  13'd173,  13'd670,  
13'd809,  13'd254,  -13'd504,  -13'd80,  -13'd812,  -13'd240,  -13'd455,  13'd348,  -13'd191,  -13'd234,  13'd75,  -13'd102,  13'd346,  13'd271,  13'd36,  13'd314,  
13'd11,  13'd529,  13'd1034,  -13'd710,  13'd122,  -13'd159,  13'd248,  -13'd2,  -13'd149,  -13'd909,  -13'd164,  -13'd108,  -13'd134,  -13'd211,  -13'd321,  13'd221,  

-13'd243,  -13'd910,  -13'd236,  13'd439,  13'd849,  -13'd252,  -13'd935,  -13'd341,  13'd11,  13'd566,  -13'd744,  13'd459,  13'd240,  -13'd846,  13'd329,  -13'd545,  
13'd617,  -13'd725,  -13'd248,  -13'd168,  13'd793,  13'd24,  -13'd224,  13'd39,  -13'd384,  13'd75,  -13'd301,  -13'd72,  13'd263,  13'd306,  13'd329,  -13'd388,  
13'd391,  -13'd82,  13'd787,  13'd212,  -13'd411,  -13'd110,  -13'd94,  13'd7,  13'd165,  -13'd312,  -13'd439,  13'd845,  -13'd555,  13'd106,  13'd498,  -13'd353,  
13'd231,  13'd60,  13'd530,  13'd481,  -13'd172,  13'd143,  13'd229,  13'd583,  -13'd335,  -13'd441,  -13'd57,  13'd205,  -13'd194,  13'd0,  13'd428,  -13'd279,  
13'd668,  13'd104,  13'd282,  13'd1093,  -13'd57,  13'd85,  -13'd51,  -13'd396,  13'd688,  -13'd137,  -13'd219,  13'd266,  -13'd41,  -13'd968,  13'd815,  -13'd449,  
-13'd67,  13'd77,  13'd334,  13'd921,  -13'd607,  13'd655,  13'd117,  -13'd265,  -13'd108,  13'd1,  -13'd459,  13'd640,  -13'd442,  13'd483,  13'd34,  -13'd81,  
13'd446,  -13'd926,  -13'd682,  13'd105,  -13'd435,  13'd467,  13'd71,  13'd421,  13'd384,  13'd338,  13'd64,  13'd29,  -13'd160,  -13'd277,  13'd345,  13'd523,  
-13'd275,  -13'd334,  -13'd146,  13'd530,  -13'd90,  -13'd328,  13'd26,  13'd59,  -13'd410,  13'd29,  -13'd571,  -13'd50,  -13'd389,  13'd1102,  13'd87,  -13'd151,  
13'd125,  13'd88,  -13'd97,  -13'd289,  -13'd83,  -13'd107,  -13'd374,  13'd965,  -13'd1003,  -13'd666,  -13'd502,  13'd209,  13'd38,  13'd180,  13'd965,  -13'd173,  
13'd905,  13'd1183,  13'd902,  -13'd353,  -13'd626,  -13'd48,  13'd139,  -13'd404,  13'd126,  -13'd996,  -13'd349,  13'd91,  -13'd896,  -13'd6,  13'd931,  13'd213,  
-13'd347,  13'd577,  13'd584,  13'd136,  13'd147,  -13'd31,  13'd1009,  -13'd124,  13'd672,  13'd269,  -13'd317,  -13'd467,  -13'd148,  -13'd156,  13'd359,  13'd242,  
13'd54,  -13'd875,  -13'd313,  -13'd483,  13'd648,  -13'd373,  13'd981,  -13'd263,  -13'd21,  -13'd482,  -13'd156,  13'd478,  13'd595,  13'd768,  13'd82,  13'd68,  
-13'd739,  13'd512,  13'd209,  -13'd321,  -13'd324,  -13'd672,  -13'd364,  13'd929,  -13'd1081,  13'd341,  -13'd53,  -13'd332,  -13'd425,  13'd252,  13'd272,  -13'd30,  
-13'd237,  -13'd34,  13'd853,  -13'd433,  -13'd640,  13'd43,  -13'd364,  13'd842,  13'd119,  -13'd870,  -13'd45,  13'd252,  -13'd988,  13'd91,  13'd808,  -13'd104,  
13'd109,  -13'd8,  13'd910,  13'd121,  -13'd540,  -13'd441,  -13'd382,  13'd523,  13'd89,  -13'd607,  -13'd703,  13'd318,  -13'd571,  -13'd307,  13'd188,  -13'd222,  
13'd7,  13'd97,  -13'd326,  -13'd50,  -13'd112,  13'd565,  13'd943,  13'd268,  -13'd627,  -13'd121,  -13'd100,  -13'd414,  13'd109,  -13'd179,  13'd339,  13'd602,  
13'd282,  -13'd39,  13'd79,  13'd748,  13'd590,  -13'd132,  -13'd168,  13'd475,  -13'd329,  -13'd521,  -13'd422,  -13'd410,  13'd184,  -13'd701,  13'd176,  -13'd559,  
-13'd559,  13'd74,  -13'd114,  -13'd424,  -13'd160,  -13'd876,  -13'd419,  13'd444,  -13'd702,  13'd498,  -13'd18,  -13'd873,  13'd115,  13'd568,  13'd8,  -13'd764,  
13'd36,  13'd25,  13'd766,  13'd83,  13'd373,  13'd466,  13'd567,  -13'd327,  13'd232,  -13'd575,  13'd182,  13'd682,  13'd128,  -13'd343,  -13'd414,  -13'd246,  
13'd1131,  13'd134,  13'd681,  -13'd58,  -13'd685,  13'd628,  13'd274,  13'd429,  -13'd671,  -13'd221,  -13'd495,  -13'd68,  13'd130,  -13'd565,  -13'd113,  13'd561,  
13'd680,  13'd446,  13'd497,  13'd293,  13'd220,  13'd427,  -13'd351,  13'd853,  -13'd516,  13'd265,  13'd78,  -13'd386,  13'd356,  13'd763,  13'd378,  -13'd41,  
-13'd394,  13'd59,  13'd894,  13'd195,  13'd49,  13'd216,  -13'd48,  13'd149,  13'd168,  13'd385,  -13'd398,  13'd282,  13'd91,  13'd598,  -13'd110,  -13'd538,  
-13'd696,  -13'd657,  -13'd64,  13'd81,  -13'd517,  -13'd184,  13'd634,  -13'd15,  -13'd523,  -13'd669,  -13'd211,  13'd177,  13'd49,  -13'd134,  13'd528,  13'd109,  
-13'd101,  13'd198,  -13'd17,  -13'd79,  13'd389,  -13'd745,  13'd253,  -13'd387,  -13'd200,  13'd1003,  13'd338,  -13'd333,  -13'd319,  -13'd302,  -13'd359,  -13'd331,  
13'd380,  13'd218,  -13'd205,  13'd69,  13'd380,  -13'd350,  13'd164,  13'd793,  -13'd509,  -13'd516,  -13'd125,  13'd277,  -13'd372,  13'd450,  -13'd542,  13'd83,  

-13'd190,  13'd181,  -13'd539,  -13'd411,  13'd375,  13'd148,  13'd291,  -13'd59,  -13'd164,  13'd167,  13'd324,  13'd306,  -13'd108,  13'd636,  -13'd356,  -13'd283,  
13'd551,  -13'd251,  13'd37,  -13'd232,  -13'd462,  13'd26,  -13'd477,  -13'd147,  13'd487,  -13'd543,  -13'd389,  -13'd79,  -13'd0,  -13'd222,  -13'd662,  13'd4,  
13'd9,  -13'd152,  -13'd586,  -13'd147,  -13'd325,  13'd76,  -13'd757,  13'd70,  -13'd501,  13'd212,  -13'd479,  -13'd86,  13'd489,  -13'd887,  -13'd51,  13'd471,  
-13'd78,  13'd40,  -13'd502,  -13'd364,  -13'd269,  -13'd187,  13'd340,  -13'd237,  -13'd202,  -13'd803,  13'd155,  -13'd692,  13'd309,  -13'd563,  -13'd128,  -13'd397,  
-13'd889,  13'd179,  -13'd582,  13'd58,  13'd81,  13'd111,  13'd407,  13'd338,  13'd207,  13'd280,  -13'd178,  13'd189,  -13'd325,  -13'd695,  13'd458,  -13'd148,  
-13'd638,  -13'd388,  -13'd404,  -13'd452,  -13'd212,  13'd698,  13'd487,  -13'd17,  -13'd347,  13'd203,  -13'd27,  13'd36,  -13'd520,  13'd70,  -13'd623,  13'd435,  
13'd216,  -13'd698,  -13'd42,  -13'd219,  -13'd596,  -13'd314,  -13'd111,  13'd341,  -13'd17,  -13'd645,  -13'd473,  -13'd193,  -13'd254,  -13'd451,  13'd128,  13'd149,  
13'd248,  13'd538,  -13'd170,  -13'd251,  13'd559,  -13'd157,  -13'd72,  -13'd714,  13'd52,  -13'd61,  13'd113,  13'd79,  -13'd423,  -13'd52,  -13'd176,  -13'd224,  
-13'd229,  -13'd544,  -13'd817,  -13'd346,  -13'd601,  13'd654,  13'd106,  -13'd415,  13'd105,  13'd318,  -13'd4,  -13'd35,  -13'd917,  -13'd607,  -13'd557,  13'd338,  
13'd163,  -13'd424,  -13'd62,  -13'd539,  -13'd279,  13'd488,  -13'd77,  13'd100,  13'd335,  13'd502,  -13'd105,  -13'd27,  13'd272,  -13'd41,  -13'd132,  13'd403,  
-13'd130,  -13'd223,  13'd232,  13'd484,  13'd15,  -13'd430,  -13'd120,  -13'd32,  -13'd836,  13'd334,  -13'd121,  -13'd327,  -13'd157,  13'd139,  13'd327,  13'd147,  
-13'd404,  -13'd315,  -13'd147,  13'd170,  -13'd193,  13'd347,  13'd21,  -13'd794,  13'd104,  13'd246,  -13'd276,  13'd602,  -13'd271,  13'd473,  -13'd102,  13'd123,  
13'd82,  -13'd67,  13'd199,  -13'd126,  13'd4,  -13'd690,  -13'd196,  -13'd371,  -13'd115,  -13'd152,  -13'd125,  13'd113,  -13'd87,  -13'd534,  13'd50,  13'd431,  
13'd297,  -13'd414,  13'd110,  13'd295,  13'd417,  13'd56,  -13'd468,  -13'd198,  -13'd53,  -13'd300,  -13'd488,  -13'd65,  -13'd607,  13'd611,  13'd365,  -13'd246,  
13'd179,  -13'd49,  -13'd445,  -13'd496,  -13'd489,  -13'd414,  13'd199,  -13'd358,  13'd515,  -13'd385,  13'd322,  -13'd336,  13'd49,  13'd38,  13'd522,  13'd270,  
-13'd147,  -13'd206,  -13'd742,  13'd217,  -13'd87,  -13'd405,  -13'd868,  13'd223,  -13'd281,  13'd241,  -13'd734,  -13'd374,  -13'd346,  13'd284,  -13'd524,  -13'd150,  
-13'd280,  -13'd378,  13'd463,  13'd91,  -13'd226,  13'd115,  -13'd24,  -13'd156,  13'd93,  13'd145,  -13'd776,  13'd9,  -13'd455,  -13'd561,  13'd306,  -13'd478,  
-13'd313,  -13'd442,  -13'd538,  13'd233,  -13'd629,  13'd59,  -13'd187,  13'd423,  -13'd554,  -13'd281,  -13'd360,  13'd61,  -13'd530,  13'd157,  -13'd673,  13'd318,  
13'd312,  13'd142,  -13'd104,  13'd159,  -13'd10,  -13'd110,  13'd300,  -13'd279,  -13'd446,  -13'd238,  -13'd20,  -13'd223,  13'd340,  -13'd351,  -13'd414,  13'd56,  
13'd129,  13'd227,  -13'd100,  13'd346,  -13'd395,  -13'd5,  -13'd725,  -13'd57,  -13'd787,  13'd336,  -13'd451,  -13'd186,  13'd273,  -13'd307,  13'd746,  13'd655,  
13'd494,  -13'd350,  13'd143,  -13'd426,  -13'd345,  -13'd110,  13'd329,  -13'd401,  -13'd293,  -13'd360,  13'd514,  13'd574,  -13'd310,  -13'd651,  -13'd616,  13'd193,  
-13'd171,  13'd532,  -13'd316,  -13'd221,  -13'd190,  13'd89,  -13'd473,  -13'd20,  -13'd423,  13'd287,  -13'd76,  13'd10,  -13'd169,  -13'd786,  -13'd482,  -13'd734,  
13'd615,  -13'd38,  13'd554,  -13'd404,  -13'd196,  13'd188,  -13'd230,  -13'd475,  -13'd269,  -13'd25,  -13'd549,  -13'd292,  -13'd61,  13'd38,  -13'd27,  13'd96,  
-13'd416,  13'd202,  -13'd154,  13'd711,  -13'd744,  -13'd439,  -13'd190,  13'd216,  13'd446,  -13'd34,  -13'd310,  -13'd679,  13'd45,  -13'd535,  13'd555,  13'd258,  
13'd399,  13'd618,  13'd259,  13'd127,  -13'd382,  -13'd178,  -13'd282,  13'd138,  -13'd390,  -13'd3,  -13'd107,  -13'd336,  13'd466,  13'd277,  13'd448,  -13'd195,  

-13'd480,  -13'd695,  -13'd627,  -13'd223,  -13'd47,  -13'd231,  -13'd1014,  13'd381,  13'd447,  13'd849,  13'd335,  -13'd53,  13'd579,  13'd298,  13'd414,  -13'd38,  
-13'd563,  13'd472,  13'd78,  13'd480,  -13'd261,  -13'd164,  -13'd676,  13'd587,  13'd24,  13'd491,  -13'd185,  -13'd10,  13'd290,  -13'd409,  13'd686,  -13'd387,  
-13'd334,  13'd320,  13'd570,  13'd833,  -13'd455,  13'd413,  -13'd34,  13'd237,  -13'd240,  -13'd715,  -13'd587,  13'd410,  13'd666,  -13'd1050,  13'd643,  13'd410,  
-13'd209,  -13'd479,  13'd97,  13'd455,  13'd128,  -13'd309,  -13'd799,  13'd596,  -13'd330,  13'd740,  13'd164,  13'd118,  -13'd550,  -13'd1425,  13'd1097,  -13'd123,  
13'd439,  -13'd243,  13'd217,  13'd190,  -13'd154,  13'd402,  13'd285,  13'd443,  13'd598,  13'd646,  13'd260,  13'd69,  -13'd69,  -13'd165,  13'd221,  -13'd410,  
13'd240,  13'd691,  13'd580,  13'd156,  -13'd491,  13'd888,  -13'd28,  -13'd4,  13'd285,  -13'd511,  -13'd381,  13'd240,  13'd597,  -13'd43,  13'd72,  -13'd174,  
13'd614,  -13'd384,  13'd9,  -13'd160,  13'd23,  -13'd49,  -13'd311,  13'd310,  13'd397,  -13'd816,  -13'd209,  13'd463,  13'd298,  13'd716,  -13'd124,  13'd432,  
-13'd189,  13'd589,  13'd6,  -13'd616,  -13'd365,  13'd806,  13'd9,  -13'd163,  -13'd36,  -13'd315,  -13'd456,  -13'd301,  -13'd417,  13'd140,  13'd138,  13'd155,  
-13'd306,  13'd629,  13'd103,  -13'd149,  -13'd335,  13'd72,  -13'd477,  13'd174,  -13'd75,  13'd506,  -13'd65,  -13'd493,  -13'd254,  13'd506,  13'd357,  13'd525,  
-13'd472,  -13'd360,  -13'd356,  13'd183,  13'd268,  -13'd393,  13'd332,  -13'd381,  -13'd387,  13'd52,  -13'd44,  13'd179,  -13'd454,  -13'd632,  13'd345,  13'd483,  
13'd461,  -13'd126,  -13'd227,  13'd342,  13'd17,  13'd44,  -13'd389,  13'd539,  13'd732,  13'd305,  -13'd1155,  -13'd134,  -13'd28,  13'd236,  13'd419,  -13'd52,  
13'd531,  -13'd217,  -13'd328,  -13'd666,  13'd256,  13'd428,  13'd489,  13'd104,  13'd331,  -13'd695,  -13'd406,  13'd88,  13'd816,  13'd195,  13'd455,  13'd541,  
-13'd479,  13'd864,  -13'd499,  -13'd725,  13'd260,  -13'd194,  13'd577,  -13'd152,  13'd199,  13'd461,  13'd224,  -13'd396,  13'd167,  13'd693,  -13'd140,  13'd200,  
13'd146,  13'd222,  13'd561,  13'd422,  -13'd37,  -13'd228,  -13'd49,  13'd144,  -13'd565,  -13'd358,  13'd101,  13'd164,  -13'd240,  13'd675,  13'd342,  13'd269,  
13'd93,  -13'd131,  13'd1165,  -13'd388,  -13'd360,  13'd380,  13'd522,  -13'd584,  -13'd450,  -13'd351,  -13'd213,  13'd241,  -13'd781,  -13'd474,  13'd294,  13'd507,  
13'd137,  13'd161,  -13'd209,  13'd45,  13'd463,  13'd219,  13'd5,  -13'd343,  -13'd521,  13'd355,  -13'd1059,  -13'd184,  13'd244,  13'd192,  -13'd91,  -13'd286,  
13'd121,  13'd356,  13'd238,  13'd179,  13'd686,  -13'd32,  13'd253,  13'd528,  -13'd26,  13'd194,  13'd557,  -13'd503,  13'd377,  -13'd491,  -13'd172,  13'd58,  
-13'd445,  13'd505,  -13'd199,  -13'd153,  -13'd443,  13'd267,  -13'd212,  -13'd264,  13'd377,  -13'd74,  -13'd470,  -13'd127,  -13'd178,  -13'd217,  -13'd167,  13'd167,  
13'd921,  13'd399,  13'd420,  13'd168,  13'd189,  13'd742,  -13'd33,  13'd28,  13'd535,  -13'd399,  13'd532,  13'd840,  13'd265,  -13'd451,  -13'd345,  -13'd138,  
13'd262,  13'd690,  -13'd159,  13'd27,  -13'd244,  -13'd106,  13'd253,  13'd195,  -13'd244,  -13'd31,  13'd40,  -13'd298,  13'd932,  -13'd233,  -13'd284,  13'd132,  
-13'd420,  13'd411,  -13'd289,  -13'd272,  -13'd151,  -13'd100,  -13'd502,  -13'd100,  -13'd47,  -13'd233,  -13'd247,  13'd462,  -13'd448,  -13'd270,  -13'd567,  -13'd107,  
-13'd18,  13'd68,  -13'd266,  13'd439,  13'd124,  13'd41,  13'd428,  -13'd344,  13'd11,  -13'd227,  13'd196,  13'd655,  -13'd502,  -13'd512,  -13'd224,  13'd762,  
-13'd722,  -13'd836,  13'd28,  -13'd578,  -13'd196,  -13'd77,  13'd331,  -13'd377,  -13'd619,  13'd367,  -13'd456,  13'd378,  13'd25,  -13'd311,  13'd108,  -13'd434,  
13'd680,  -13'd439,  13'd327,  -13'd238,  -13'd82,  -13'd374,  13'd338,  -13'd182,  -13'd243,  13'd377,  13'd132,  -13'd717,  13'd202,  13'd1061,  -13'd941,  13'd388,  
-13'd492,  -13'd600,  -13'd165,  -13'd341,  13'd78,  -13'd270,  13'd343,  -13'd331,  -13'd214,  -13'd1199,  -13'd948,  -13'd352,  13'd259,  -13'd334,  -13'd838,  13'd268,  

13'd325,  13'd233,  -13'd456,  13'd415,  13'd347,  13'd178,  13'd228,  -13'd186,  13'd138,  -13'd699,  13'd1509,  13'd169,  -13'd282,  -13'd373,  -13'd374,  -13'd933,  
-13'd736,  -13'd550,  -13'd670,  13'd365,  -13'd630,  -13'd460,  -13'd1046,  -13'd681,  13'd357,  -13'd291,  13'd558,  13'd216,  -13'd546,  -13'd402,  -13'd553,  -13'd457,  
13'd199,  13'd223,  -13'd219,  13'd437,  -13'd44,  13'd810,  -13'd885,  13'd738,  13'd147,  13'd125,  13'd62,  -13'd30,  -13'd443,  -13'd1418,  -13'd430,  13'd684,  
-13'd865,  -13'd624,  13'd505,  -13'd663,  -13'd500,  13'd5,  -13'd44,  -13'd304,  13'd856,  13'd709,  13'd125,  -13'd341,  13'd403,  -13'd1026,  -13'd65,  13'd144,  
-13'd216,  -13'd939,  13'd843,  -13'd109,  -13'd99,  -13'd707,  -13'd34,  13'd133,  13'd183,  13'd437,  13'd189,  -13'd406,  -13'd626,  -13'd181,  -13'd1022,  13'd97,  
13'd529,  13'd22,  13'd273,  13'd669,  13'd160,  13'd517,  -13'd717,  13'd130,  13'd703,  13'd513,  13'd234,  13'd222,  13'd227,  -13'd80,  13'd49,  13'd68,  
13'd100,  13'd462,  13'd164,  -13'd208,  -13'd499,  13'd18,  -13'd340,  -13'd262,  13'd111,  -13'd65,  -13'd271,  -13'd212,  13'd88,  13'd22,  13'd212,  13'd607,  
13'd56,  -13'd348,  -13'd60,  13'd796,  -13'd380,  13'd182,  -13'd798,  13'd22,  -13'd162,  13'd322,  -13'd236,  13'd164,  -13'd440,  -13'd561,  13'd476,  13'd88,  
-13'd712,  13'd152,  -13'd407,  -13'd68,  -13'd342,  -13'd160,  13'd670,  -13'd345,  13'd504,  13'd552,  -13'd504,  -13'd703,  13'd166,  13'd87,  -13'd124,  -13'd226,  
-13'd650,  -13'd164,  -13'd467,  13'd537,  -13'd77,  -13'd126,  -13'd374,  13'd526,  -13'd54,  13'd582,  -13'd105,  -13'd184,  13'd64,  -13'd371,  -13'd859,  -13'd300,  
13'd177,  -13'd140,  -13'd15,  13'd255,  13'd666,  13'd240,  13'd108,  13'd565,  -13'd7,  13'd53,  13'd53,  -13'd317,  13'd305,  13'd196,  13'd436,  -13'd85,  
-13'd591,  13'd175,  -13'd10,  13'd724,  13'd580,  -13'd707,  -13'd159,  -13'd489,  13'd785,  -13'd348,  13'd881,  13'd5,  13'd277,  -13'd333,  13'd167,  13'd192,  
13'd280,  13'd453,  -13'd245,  13'd208,  -13'd102,  -13'd412,  -13'd15,  13'd528,  -13'd523,  -13'd61,  13'd625,  13'd230,  -13'd104,  -13'd513,  -13'd4,  13'd233,  
13'd843,  -13'd53,  13'd99,  -13'd505,  13'd147,  -13'd22,  13'd591,  13'd341,  -13'd333,  -13'd909,  13'd565,  -13'd148,  13'd143,  -13'd495,  13'd355,  13'd173,  
-13'd217,  13'd421,  13'd320,  -13'd137,  13'd595,  13'd662,  13'd306,  -13'd146,  -13'd135,  13'd376,  13'd240,  -13'd96,  13'd601,  13'd38,  -13'd395,  -13'd321,  
-13'd496,  13'd707,  13'd453,  13'd541,  13'd1008,  -13'd321,  -13'd781,  13'd178,  -13'd24,  13'd119,  -13'd279,  -13'd268,  13'd306,  13'd9,  -13'd121,  13'd49,  
-13'd410,  13'd386,  -13'd208,  13'd455,  13'd597,  -13'd221,  -13'd1009,  13'd269,  13'd635,  -13'd743,  13'd138,  -13'd229,  13'd321,  -13'd1026,  13'd288,  -13'd11,  
13'd605,  -13'd604,  13'd577,  -13'd500,  -13'd524,  -13'd613,  -13'd336,  13'd17,  -13'd43,  -13'd37,  -13'd575,  13'd746,  -13'd285,  13'd909,  -13'd559,  -13'd251,  
13'd836,  13'd63,  13'd634,  -13'd419,  -13'd672,  -13'd219,  13'd681,  -13'd535,  13'd395,  -13'd172,  13'd190,  13'd713,  13'd416,  13'd149,  13'd164,  13'd256,  
-13'd184,  -13'd228,  -13'd951,  -13'd168,  -13'd188,  -13'd210,  -13'd384,  13'd646,  -13'd427,  13'd109,  13'd429,  13'd34,  -13'd196,  13'd64,  13'd596,  13'd534,  
-13'd687,  13'd964,  -13'd435,  -13'd710,  13'd150,  -13'd721,  13'd1009,  -13'd539,  13'd523,  -13'd51,  -13'd519,  13'd121,  13'd251,  -13'd493,  -13'd125,  -13'd157,  
-13'd38,  -13'd175,  -13'd487,  -13'd339,  -13'd189,  13'd214,  13'd1067,  13'd290,  13'd368,  -13'd753,  13'd263,  13'd201,  -13'd34,  -13'd461,  -13'd390,  -13'd583,  
-13'd683,  -13'd81,  -13'd124,  13'd84,  -13'd582,  -13'd484,  13'd491,  -13'd819,  13'd783,  13'd333,  13'd514,  -13'd50,  -13'd212,  13'd658,  13'd540,  13'd464,  
-13'd585,  -13'd381,  -13'd204,  13'd690,  13'd711,  -13'd477,  13'd490,  -13'd472,  -13'd88,  13'd168,  -13'd454,  13'd127,  -13'd114,  -13'd370,  13'd111,  -13'd148,  
-13'd505,  -13'd355,  13'd533,  -13'd67,  -13'd568,  13'd441,  13'd53,  -13'd183,  -13'd101,  13'd876,  -13'd562,  13'd535,  -13'd69,  13'd158,  13'd372,  13'd260,  

13'd326,  -13'd307,  13'd600,  -13'd500,  -13'd767,  -13'd386,  13'd197,  13'd1,  -13'd132,  13'd417,  13'd721,  -13'd338,  -13'd285,  -13'd65,  -13'd19,  -13'd349,  
-13'd613,  -13'd445,  -13'd1064,  -13'd278,  -13'd173,  13'd146,  13'd296,  13'd353,  13'd531,  -13'd587,  13'd307,  13'd771,  13'd591,  -13'd658,  -13'd106,  -13'd83,  
13'd43,  13'd83,  -13'd763,  13'd400,  13'd868,  13'd513,  13'd44,  13'd241,  -13'd559,  13'd289,  13'd868,  13'd397,  13'd267,  -13'd418,  -13'd471,  -13'd290,  
13'd878,  13'd718,  13'd287,  13'd710,  -13'd60,  13'd353,  -13'd96,  13'd35,  13'd321,  13'd439,  13'd203,  -13'd46,  -13'd227,  -13'd1098,  13'd26,  13'd432,  
-13'd32,  13'd286,  13'd13,  -13'd243,  13'd406,  13'd463,  13'd399,  13'd804,  -13'd307,  -13'd181,  13'd91,  -13'd347,  13'd1012,  -13'd327,  -13'd658,  -13'd505,  
-13'd393,  -13'd758,  13'd317,  -13'd472,  13'd144,  -13'd72,  -13'd676,  -13'd191,  13'd777,  13'd333,  13'd416,  13'd474,  13'd45,  -13'd479,  13'd483,  -13'd745,  
13'd507,  13'd390,  13'd279,  -13'd735,  -13'd37,  -13'd754,  13'd306,  -13'd792,  -13'd622,  -13'd311,  13'd96,  -13'd130,  13'd260,  -13'd372,  -13'd397,  13'd141,  
-13'd430,  13'd65,  13'd293,  13'd426,  13'd514,  13'd420,  13'd826,  -13'd403,  -13'd653,  13'd99,  13'd484,  13'd459,  -13'd78,  -13'd736,  13'd705,  -13'd464,  
13'd421,  13'd190,  -13'd951,  13'd208,  13'd900,  13'd115,  13'd132,  13'd32,  13'd80,  -13'd360,  13'd475,  -13'd469,  13'd399,  -13'd451,  13'd532,  13'd220,  
-13'd1601,  -13'd109,  -13'd1010,  13'd362,  -13'd255,  -13'd528,  13'd24,  -13'd428,  13'd535,  13'd793,  13'd476,  13'd130,  13'd633,  13'd343,  -13'd23,  13'd889,  
13'd359,  -13'd83,  13'd242,  13'd525,  -13'd198,  -13'd57,  13'd643,  -13'd528,  -13'd493,  -13'd239,  -13'd749,  -13'd155,  -13'd184,  13'd180,  13'd645,  13'd482,  
13'd673,  -13'd270,  13'd247,  13'd587,  -13'd777,  13'd165,  13'd295,  -13'd164,  -13'd161,  -13'd808,  13'd900,  13'd161,  13'd288,  -13'd529,  13'd74,  -13'd576,  
13'd148,  -13'd715,  -13'd188,  13'd60,  -13'd271,  -13'd29,  13'd711,  13'd348,  13'd578,  13'd211,  13'd942,  -13'd487,  13'd636,  -13'd497,  13'd36,  -13'd100,  
13'd106,  13'd23,  -13'd253,  13'd212,  -13'd661,  13'd56,  -13'd514,  -13'd238,  13'd501,  -13'd556,  13'd260,  13'd126,  13'd91,  -13'd23,  13'd554,  13'd84,  
-13'd1096,  -13'd492,  -13'd91,  13'd727,  -13'd206,  13'd150,  -13'd86,  -13'd119,  13'd203,  13'd1534,  13'd771,  13'd601,  -13'd680,  13'd709,  -13'd72,  -13'd994,  
13'd28,  13'd282,  -13'd1,  13'd733,  -13'd109,  13'd260,  -13'd238,  -13'd137,  13'd370,  13'd520,  13'd463,  13'd648,  -13'd38,  -13'd477,  -13'd609,  13'd832,  
13'd837,  -13'd624,  13'd321,  13'd780,  -13'd230,  13'd341,  13'd1267,  13'd742,  -13'd130,  -13'd816,  13'd257,  13'd53,  13'd696,  -13'd252,  13'd32,  13'd443,  
-13'd475,  13'd566,  -13'd143,  -13'd378,  -13'd234,  13'd206,  13'd285,  -13'd37,  13'd143,  -13'd90,  -13'd503,  13'd381,  -13'd280,  -13'd248,  -13'd215,  -13'd224,  
13'd588,  13'd84,  13'd691,  -13'd450,  -13'd1021,  -13'd234,  13'd235,  13'd834,  13'd698,  13'd132,  13'd133,  -13'd289,  -13'd238,  -13'd205,  13'd79,  13'd428,  
13'd606,  -13'd177,  -13'd984,  13'd469,  13'd77,  -13'd686,  13'd164,  13'd509,  13'd796,  13'd208,  13'd227,  13'd296,  -13'd522,  13'd571,  13'd199,  -13'd157,  
13'd603,  13'd345,  -13'd36,  -13'd1234,  -13'd507,  13'd232,  13'd361,  -13'd34,  -13'd1051,  -13'd164,  13'd411,  13'd366,  -13'd520,  13'd35,  -13'd686,  13'd226,  
13'd317,  -13'd213,  13'd1295,  -13'd136,  -13'd57,  -13'd136,  13'd845,  -13'd652,  13'd275,  13'd141,  -13'd414,  -13'd681,  13'd130,  13'd131,  -13'd438,  13'd671,  
-13'd201,  13'd341,  13'd124,  -13'd765,  13'd883,  -13'd254,  13'd514,  13'd83,  13'd1195,  -13'd85,  -13'd639,  -13'd1050,  -13'd602,  13'd1162,  13'd532,  -13'd633,  
-13'd109,  -13'd1003,  13'd223,  13'd162,  -13'd226,  -13'd625,  -13'd566,  -13'd892,  13'd988,  -13'd4,  -13'd717,  -13'd786,  -13'd1095,  -13'd158,  -13'd84,  -13'd570,  
-13'd244,  -13'd881,  13'd13,  13'd28,  -13'd49,  13'd1114,  13'd16,  -13'd184,  13'd394,  13'd978,  -13'd473,  -13'd305,  -13'd297,  13'd200,  13'd464,  -13'd67,  

13'd116,  -13'd741,  -13'd73,  -13'd91,  -13'd112,  13'd175,  -13'd270,  13'd674,  13'd887,  -13'd163,  -13'd168,  13'd248,  13'd306,  13'd198,  -13'd587,  -13'd120,  
13'd193,  13'd310,  13'd222,  -13'd673,  13'd346,  -13'd14,  13'd47,  13'd581,  13'd647,  -13'd53,  13'd552,  -13'd71,  -13'd17,  -13'd703,  13'd295,  -13'd432,  
13'd8,  -13'd292,  -13'd124,  13'd250,  13'd134,  13'd328,  -13'd400,  13'd11,  -13'd470,  13'd126,  -13'd202,  -13'd7,  -13'd79,  -13'd177,  13'd49,  -13'd203,  
-13'd64,  -13'd182,  -13'd159,  -13'd186,  -13'd73,  -13'd577,  13'd309,  13'd307,  13'd146,  -13'd22,  -13'd57,  -13'd12,  -13'd620,  -13'd78,  -13'd313,  -13'd137,  
-13'd179,  -13'd624,  13'd715,  -13'd303,  -13'd229,  -13'd22,  -13'd729,  -13'd60,  13'd468,  13'd137,  -13'd188,  13'd261,  -13'd59,  -13'd672,  13'd243,  -13'd38,  
-13'd334,  13'd473,  13'd214,  13'd107,  13'd16,  13'd398,  -13'd434,  -13'd39,  13'd469,  -13'd272,  -13'd290,  -13'd30,  13'd327,  -13'd728,  13'd556,  13'd71,  
-13'd172,  13'd111,  13'd0,  -13'd8,  -13'd202,  13'd430,  13'd372,  13'd241,  -13'd162,  -13'd476,  -13'd155,  -13'd388,  -13'd427,  13'd5,  -13'd585,  13'd566,  
13'd50,  -13'd378,  13'd619,  13'd432,  13'd214,  -13'd52,  -13'd702,  -13'd139,  -13'd683,  -13'd123,  -13'd158,  -13'd511,  13'd146,  -13'd449,  13'd332,  -13'd272,  
-13'd413,  -13'd428,  -13'd722,  13'd160,  -13'd81,  13'd9,  -13'd574,  13'd210,  -13'd67,  -13'd660,  13'd30,  -13'd97,  -13'd401,  -13'd146,  -13'd572,  -13'd530,  
-13'd53,  -13'd324,  13'd402,  13'd110,  13'd192,  -13'd168,  13'd0,  -13'd6,  -13'd703,  -13'd672,  13'd496,  -13'd203,  -13'd161,  13'd697,  13'd95,  -13'd316,  
-13'd19,  13'd40,  -13'd649,  -13'd161,  13'd307,  13'd245,  13'd232,  13'd194,  -13'd284,  13'd657,  13'd275,  -13'd470,  13'd191,  -13'd358,  -13'd105,  -13'd250,  
-13'd451,  13'd664,  -13'd438,  13'd401,  -13'd465,  13'd6,  -13'd248,  13'd133,  13'd128,  -13'd450,  -13'd375,  13'd350,  -13'd334,  13'd249,  -13'd874,  -13'd222,  
-13'd369,  -13'd57,  13'd71,  13'd402,  -13'd140,  13'd766,  -13'd603,  -13'd355,  -13'd433,  -13'd331,  -13'd8,  13'd271,  13'd96,  -13'd287,  13'd418,  -13'd483,  
13'd10,  13'd207,  -13'd488,  -13'd210,  13'd323,  -13'd330,  -13'd8,  -13'd596,  -13'd669,  -13'd595,  -13'd467,  -13'd654,  -13'd176,  13'd58,  13'd131,  -13'd329,  
13'd445,  13'd120,  13'd526,  13'd717,  -13'd587,  -13'd37,  13'd372,  -13'd290,  -13'd122,  13'd134,  -13'd219,  -13'd282,  13'd264,  -13'd122,  13'd163,  -13'd727,  
13'd474,  13'd184,  13'd169,  -13'd422,  13'd212,  13'd459,  13'd15,  13'd2,  13'd300,  13'd347,  -13'd209,  -13'd212,  -13'd391,  -13'd470,  -13'd701,  13'd3,  
13'd7,  -13'd444,  13'd222,  13'd87,  13'd297,  -13'd808,  -13'd548,  13'd243,  13'd157,  -13'd6,  13'd298,  -13'd82,  -13'd159,  -13'd478,  -13'd165,  -13'd417,  
13'd25,  -13'd270,  13'd2,  -13'd306,  13'd78,  -13'd207,  -13'd449,  -13'd642,  -13'd391,  13'd341,  13'd290,  -13'd230,  13'd197,  13'd658,  13'd117,  -13'd460,  
13'd9,  13'd466,  -13'd304,  -13'd589,  -13'd713,  -13'd585,  -13'd415,  -13'd321,  13'd160,  -13'd199,  13'd32,  -13'd514,  -13'd266,  13'd200,  -13'd249,  13'd147,  
-13'd582,  -13'd158,  -13'd66,  -13'd528,  13'd448,  13'd271,  13'd146,  -13'd251,  -13'd518,  -13'd396,  -13'd495,  -13'd577,  -13'd607,  13'd407,  -13'd81,  -13'd184,  
-13'd580,  -13'd42,  -13'd489,  13'd103,  13'd43,  13'd177,  -13'd189,  13'd221,  13'd562,  -13'd107,  13'd520,  -13'd61,  13'd269,  -13'd795,  13'd208,  13'd587,  
-13'd446,  -13'd359,  13'd673,  13'd196,  13'd17,  13'd595,  -13'd613,  -13'd197,  -13'd143,  13'd482,  -13'd406,  13'd295,  -13'd36,  -13'd171,  13'd84,  -13'd180,  
13'd147,  -13'd435,  -13'd243,  -13'd785,  13'd270,  -13'd404,  13'd295,  13'd8,  -13'd295,  13'd114,  -13'd218,  -13'd164,  13'd80,  -13'd323,  13'd95,  13'd34,  
-13'd352,  -13'd371,  13'd239,  13'd355,  -13'd540,  -13'd381,  -13'd131,  -13'd585,  -13'd265,  13'd93,  -13'd658,  -13'd656,  13'd59,  -13'd131,  -13'd120,  -13'd45,  
-13'd158,  13'd676,  13'd561,  -13'd97,  -13'd690,  13'd37,  -13'd103,  -13'd344,  -13'd285,  -13'd2,  -13'd825,  13'd445,  -13'd417,  -13'd408,  -13'd646,  -13'd26,  

-13'd392,  13'd51,  13'd834,  13'd801,  13'd25,  -13'd111,  -13'd511,  13'd717,  -13'd102,  13'd432,  13'd60,  -13'd1104,  13'd573,  13'd410,  -13'd109,  13'd78,  
-13'd655,  -13'd22,  13'd908,  13'd393,  -13'd142,  -13'd457,  13'd40,  13'd291,  13'd362,  -13'd5,  13'd128,  -13'd269,  13'd314,  13'd1864,  13'd436,  -13'd164,  
-13'd344,  -13'd185,  13'd1116,  13'd56,  -13'd1018,  -13'd42,  13'd463,  -13'd32,  -13'd128,  13'd385,  -13'd289,  13'd353,  -13'd226,  13'd1443,  13'd123,  -13'd470,  
13'd1029,  13'd275,  13'd444,  -13'd24,  13'd93,  13'd521,  13'd293,  -13'd575,  13'd790,  -13'd26,  13'd521,  13'd774,  -13'd459,  -13'd222,  -13'd34,  -13'd958,  
13'd946,  13'd1247,  -13'd908,  13'd557,  -13'd649,  13'd416,  13'd658,  13'd393,  13'd249,  -13'd421,  13'd686,  -13'd124,  13'd681,  -13'd833,  -13'd294,  13'd1013,  
-13'd103,  13'd556,  -13'd215,  -13'd660,  13'd1080,  -13'd569,  -13'd512,  -13'd327,  -13'd622,  -13'd574,  13'd439,  13'd278,  13'd388,  13'd610,  13'd403,  -13'd403,  
-13'd387,  -13'd112,  13'd845,  13'd285,  -13'd173,  13'd493,  13'd392,  -13'd730,  -13'd301,  -13'd86,  13'd56,  13'd157,  13'd66,  13'd997,  13'd14,  -13'd58,  
-13'd170,  -13'd339,  13'd841,  13'd500,  -13'd412,  13'd426,  -13'd19,  -13'd377,  13'd652,  -13'd541,  -13'd51,  -13'd491,  -13'd406,  13'd1168,  -13'd279,  -13'd641,  
13'd141,  -13'd345,  -13'd153,  13'd428,  -13'd396,  -13'd36,  13'd175,  13'd140,  -13'd80,  -13'd464,  -13'd324,  13'd184,  13'd503,  13'd245,  -13'd359,  -13'd339,  
13'd699,  -13'd401,  -13'd1179,  13'd322,  13'd165,  -13'd461,  -13'd208,  -13'd307,  13'd762,  13'd587,  13'd310,  -13'd425,  -13'd352,  -13'd750,  -13'd504,  13'd517,  
-13'd31,  -13'd539,  13'd63,  13'd337,  -13'd132,  -13'd633,  -13'd352,  13'd127,  -13'd474,  -13'd217,  13'd248,  13'd185,  -13'd251,  -13'd312,  13'd378,  -13'd127,  
-13'd257,  -13'd215,  -13'd294,  -13'd375,  -13'd26,  -13'd179,  -13'd46,  -13'd65,  -13'd542,  -13'd238,  -13'd387,  -13'd321,  -13'd547,  13'd905,  -13'd164,  13'd587,  
13'd192,  -13'd438,  13'd744,  -13'd594,  -13'd629,  13'd440,  -13'd78,  13'd163,  -13'd420,  13'd427,  -13'd777,  -13'd127,  -13'd243,  13'd452,  13'd71,  13'd128,  
13'd575,  13'd243,  13'd780,  13'd851,  -13'd632,  13'd693,  -13'd170,  -13'd318,  13'd398,  -13'd936,  13'd2,  13'd99,  -13'd508,  13'd470,  -13'd640,  -13'd6,  
-13'd311,  -13'd679,  13'd451,  13'd606,  -13'd355,  13'd128,  -13'd353,  -13'd264,  13'd441,  -13'd167,  -13'd284,  -13'd533,  -13'd965,  -13'd501,  13'd356,  13'd202,  
-13'd572,  13'd492,  -13'd605,  13'd568,  13'd594,  13'd199,  13'd765,  13'd720,  13'd663,  13'd169,  13'd454,  -13'd527,  13'd519,  -13'd705,  -13'd671,  -13'd93,  
-13'd427,  -13'd635,  13'd273,  13'd114,  -13'd941,  -13'd756,  13'd303,  13'd229,  13'd93,  13'd1005,  13'd406,  -13'd241,  13'd158,  -13'd348,  -13'd281,  13'd29,  
13'd166,  -13'd100,  -13'd268,  13'd479,  -13'd41,  13'd172,  13'd108,  13'd12,  -13'd16,  13'd273,  13'd28,  13'd51,  13'd457,  13'd872,  13'd148,  -13'd682,  
-13'd796,  -13'd95,  13'd168,  13'd650,  -13'd339,  -13'd493,  13'd319,  13'd674,  -13'd126,  -13'd488,  13'd675,  -13'd279,  13'd199,  -13'd324,  -13'd551,  13'd664,  
13'd368,  -13'd153,  13'd380,  13'd71,  13'd861,  -13'd223,  13'd173,  13'd43,  -13'd232,  -13'd302,  -13'd223,  13'd517,  13'd454,  13'd224,  13'd125,  13'd19,  
13'd19,  13'd469,  13'd196,  -13'd684,  -13'd752,  -13'd17,  13'd80,  -13'd580,  -13'd315,  13'd200,  13'd28,  13'd194,  -13'd390,  -13'd427,  13'd90,  13'd751,  
13'd242,  13'd504,  13'd939,  -13'd861,  13'd206,  13'd64,  13'd790,  -13'd216,  -13'd34,  13'd144,  13'd195,  13'd226,  13'd511,  13'd692,  13'd354,  -13'd38,  
-13'd48,  13'd283,  13'd276,  13'd248,  -13'd650,  -13'd127,  13'd321,  -13'd697,  -13'd22,  13'd31,  -13'd800,  -13'd410,  13'd669,  13'd844,  -13'd124,  13'd40,  
-13'd1016,  13'd542,  -13'd1112,  -13'd191,  13'd231,  -13'd87,  13'd256,  -13'd403,  -13'd423,  -13'd51,  13'd622,  -13'd1277,  13'd85,  -13'd559,  13'd366,  13'd340,  
-13'd792,  13'd85,  -13'd708,  13'd22,  13'd68,  -13'd95,  -13'd125,  13'd455,  -13'd821,  -13'd999,  13'd215,  -13'd1025,  -13'd610,  13'd548,  -13'd190,  -13'd138,  

-13'd968,  -13'd517,  13'd114,  -13'd395,  13'd1229,  13'd196,  -13'd609,  13'd886,  -13'd284,  -13'd140,  13'd266,  -13'd355,  13'd20,  -13'd975,  -13'd96,  13'd27,  
13'd44,  13'd793,  13'd418,  -13'd88,  13'd614,  13'd398,  -13'd84,  13'd662,  -13'd267,  13'd658,  -13'd684,  -13'd469,  13'd584,  -13'd328,  13'd211,  13'd560,  
-13'd546,  -13'd428,  13'd486,  13'd232,  -13'd551,  13'd336,  13'd49,  -13'd465,  -13'd898,  13'd94,  -13'd436,  -13'd145,  13'd243,  13'd260,  13'd477,  13'd322,  
-13'd341,  13'd688,  13'd612,  13'd171,  13'd57,  13'd333,  13'd161,  13'd158,  13'd581,  13'd227,  13'd558,  13'd306,  -13'd796,  13'd1125,  -13'd889,  13'd28,  
13'd929,  13'd792,  -13'd363,  13'd346,  -13'd3,  13'd494,  13'd509,  -13'd591,  13'd808,  -13'd235,  13'd407,  13'd125,  -13'd248,  13'd467,  13'd344,  13'd748,  
-13'd804,  -13'd59,  -13'd1197,  -13'd348,  -13'd332,  -13'd141,  13'd146,  13'd266,  -13'd338,  -13'd63,  13'd790,  -13'd646,  -13'd599,  -13'd834,  -13'd503,  13'd236,  
-13'd733,  -13'd431,  -13'd469,  -13'd329,  13'd995,  -13'd207,  -13'd582,  13'd172,  -13'd266,  13'd50,  13'd198,  -13'd326,  -13'd560,  -13'd556,  -13'd510,  -13'd48,  
13'd575,  -13'd411,  13'd674,  13'd206,  13'd437,  -13'd246,  13'd235,  -13'd19,  -13'd1091,  13'd423,  -13'd129,  13'd636,  -13'd59,  -13'd65,  -13'd320,  13'd89,  
13'd724,  -13'd112,  13'd904,  13'd279,  13'd688,  -13'd112,  13'd527,  13'd285,  13'd253,  -13'd631,  13'd368,  -13'd204,  13'd229,  13'd607,  13'd308,  -13'd218,  
13'd720,  -13'd47,  -13'd8,  13'd380,  -13'd31,  -13'd15,  13'd685,  13'd144,  13'd361,  13'd272,  -13'd211,  -13'd598,  13'd284,  -13'd302,  -13'd320,  13'd258,  
-13'd762,  -13'd505,  -13'd935,  -13'd548,  13'd398,  -13'd579,  -13'd577,  13'd277,  13'd838,  -13'd445,  13'd1119,  -13'd30,  -13'd571,  -13'd626,  13'd214,  -13'd590,  
13'd270,  13'd194,  -13'd172,  13'd262,  -13'd82,  13'd496,  -13'd493,  13'd504,  -13'd207,  13'd2,  13'd8,  -13'd138,  -13'd419,  13'd355,  13'd382,  13'd119,  
13'd922,  -13'd425,  -13'd36,  -13'd663,  13'd134,  -13'd10,  -13'd523,  13'd433,  13'd353,  13'd534,  -13'd160,  -13'd138,  13'd826,  -13'd780,  -13'd425,  13'd187,  
13'd24,  -13'd711,  -13'd140,  13'd598,  13'd485,  -13'd183,  -13'd117,  13'd619,  -13'd419,  13'd669,  13'd290,  -13'd233,  13'd753,  -13'd32,  -13'd580,  13'd325,  
-13'd897,  13'd152,  -13'd378,  13'd355,  13'd291,  -13'd621,  13'd479,  -13'd489,  -13'd500,  13'd333,  13'd228,  13'd197,  -13'd4,  -13'd543,  13'd382,  13'd338,  
13'd335,  13'd225,  -13'd582,  13'd427,  -13'd546,  -13'd112,  -13'd157,  -13'd367,  13'd474,  -13'd407,  13'd187,  -13'd110,  -13'd391,  13'd656,  -13'd34,  -13'd438,  
13'd105,  -13'd396,  -13'd47,  13'd452,  -13'd557,  13'd253,  13'd97,  13'd116,  13'd339,  13'd392,  -13'd273,  -13'd479,  13'd402,  13'd746,  13'd766,  -13'd568,  
-13'd285,  13'd83,  13'd84,  13'd338,  13'd495,  13'd71,  13'd133,  -13'd360,  -13'd185,  -13'd521,  13'd639,  13'd626,  -13'd162,  13'd126,  -13'd400,  13'd517,  
-13'd129,  -13'd24,  -13'd287,  13'd283,  13'd93,  13'd340,  13'd437,  13'd155,  13'd522,  13'd601,  13'd318,  -13'd21,  -13'd631,  -13'd420,  13'd598,  13'd374,  
13'd228,  -13'd949,  -13'd681,  13'd128,  13'd516,  -13'd265,  -13'd404,  13'd220,  -13'd336,  13'd376,  13'd1104,  13'd503,  13'd226,  13'd18,  -13'd298,  13'd758,  
13'd335,  -13'd69,  13'd730,  13'd722,  -13'd189,  -13'd86,  -13'd150,  -13'd209,  13'd436,  13'd40,  -13'd106,  -13'd27,  13'd183,  -13'd158,  13'd223,  13'd448,  
-13'd532,  -13'd284,  -13'd79,  13'd875,  13'd55,  13'd587,  -13'd524,  -13'd336,  -13'd596,  13'd506,  -13'd163,  -13'd122,  13'd162,  13'd596,  13'd610,  13'd216,  
13'd297,  13'd280,  13'd173,  -13'd43,  13'd139,  -13'd406,  -13'd515,  -13'd241,  -13'd504,  -13'd437,  -13'd105,  -13'd176,  13'd698,  -13'd267,  13'd310,  13'd648,  
-13'd52,  13'd566,  13'd224,  -13'd143,  -13'd354,  13'd27,  -13'd307,  -13'd422,  -13'd445,  -13'd604,  13'd591,  13'd49,  13'd368,  13'd247,  -13'd152,  13'd74,  
-13'd75,  13'd1023,  13'd248,  -13'd456,  13'd517,  13'd42,  -13'd372,  13'd486,  -13'd411,  -13'd223,  13'd15,  -13'd114,  -13'd225,  13'd442,  -13'd103,  13'd181,  

-13'd274,  -13'd514,  -13'd587,  -13'd353,  13'd632,  13'd159,  13'd237,  13'd522,  -13'd489,  13'd420,  13'd551,  -13'd82,  13'd1381,  -13'd199,  -13'd80,  -13'd588,  
13'd495,  -13'd190,  13'd17,  13'd433,  13'd83,  13'd435,  -13'd107,  13'd513,  -13'd456,  -13'd62,  13'd508,  13'd408,  13'd28,  13'd130,  13'd410,  13'd497,  
13'd975,  13'd267,  13'd250,  13'd371,  -13'd139,  13'd91,  -13'd304,  13'd245,  -13'd472,  -13'd717,  13'd354,  13'd23,  13'd277,  13'd202,  -13'd53,  13'd1,  
13'd68,  13'd253,  -13'd357,  13'd452,  -13'd120,  -13'd36,  -13'd2,  -13'd458,  -13'd514,  -13'd379,  13'd1116,  -13'd34,  13'd733,  -13'd148,  -13'd179,  13'd51,  
-13'd89,  -13'd600,  -13'd692,  13'd783,  13'd463,  13'd231,  -13'd216,  13'd511,  -13'd124,  -13'd555,  13'd442,  -13'd488,  13'd505,  13'd594,  -13'd38,  -13'd332,  
13'd386,  13'd395,  -13'd531,  -13'd45,  13'd645,  -13'd264,  -13'd26,  -13'd126,  -13'd446,  -13'd373,  13'd690,  -13'd533,  13'd563,  -13'd433,  13'd23,  -13'd293,  
-13'd361,  13'd185,  -13'd372,  13'd235,  -13'd56,  13'd103,  13'd125,  13'd475,  -13'd412,  -13'd274,  13'd530,  -13'd799,  -13'd252,  -13'd539,  13'd18,  -13'd49,  
-13'd186,  13'd184,  13'd514,  13'd170,  13'd555,  13'd316,  -13'd144,  13'd344,  -13'd419,  13'd18,  13'd757,  -13'd399,  13'd444,  13'd1301,  -13'd278,  13'd741,  
-13'd659,  13'd246,  13'd14,  -13'd24,  13'd55,  -13'd145,  -13'd76,  13'd565,  13'd635,  13'd291,  13'd802,  -13'd455,  -13'd97,  13'd120,  13'd410,  13'd274,  
13'd157,  13'd68,  13'd592,  -13'd114,  13'd195,  -13'd304,  13'd777,  13'd4,  13'd268,  -13'd141,  13'd917,  13'd721,  13'd89,  13'd247,  13'd112,  13'd174,  
-13'd642,  13'd904,  -13'd355,  -13'd483,  13'd303,  -13'd904,  -13'd192,  13'd141,  13'd823,  13'd154,  13'd1191,  -13'd506,  13'd61,  13'd1,  -13'd132,  -13'd416,  
-13'd502,  -13'd270,  -13'd71,  -13'd465,  13'd410,  13'd135,  -13'd646,  -13'd30,  13'd150,  13'd836,  -13'd423,  -13'd183,  -13'd914,  -13'd627,  -13'd507,  -13'd85,  
13'd113,  -13'd105,  13'd204,  -13'd707,  13'd650,  13'd176,  -13'd192,  13'd35,  13'd361,  13'd860,  13'd246,  13'd694,  13'd372,  -13'd33,  13'd286,  13'd235,  
13'd377,  13'd130,  13'd268,  13'd196,  13'd446,  13'd323,  13'd119,  -13'd145,  13'd816,  -13'd195,  13'd141,  13'd713,  -13'd203,  13'd395,  13'd728,  13'd84,  
-13'd826,  13'd68,  -13'd850,  13'd132,  -13'd161,  -13'd1161,  13'd41,  -13'd184,  13'd176,  13'd221,  -13'd29,  -13'd396,  13'd439,  13'd186,  13'd589,  -13'd312,  
13'd134,  -13'd673,  -13'd89,  -13'd49,  -13'd1008,  13'd166,  -13'd110,  -13'd149,  13'd319,  -13'd629,  -13'd224,  -13'd188,  13'd149,  -13'd186,  -13'd461,  -13'd80,  
-13'd432,  -13'd695,  -13'd525,  13'd326,  -13'd873,  13'd217,  13'd319,  13'd385,  13'd490,  13'd585,  13'd217,  13'd816,  -13'd267,  13'd521,  13'd411,  -13'd648,  
-13'd208,  -13'd49,  13'd277,  13'd156,  13'd360,  13'd426,  13'd217,  -13'd24,  -13'd54,  -13'd288,  13'd539,  13'd142,  13'd457,  -13'd499,  13'd996,  -13'd760,  
-13'd566,  -13'd367,  13'd68,  13'd100,  13'd178,  13'd326,  13'd78,  -13'd19,  13'd215,  13'd76,  -13'd241,  -13'd81,  13'd147,  -13'd430,  -13'd40,  -13'd466,  
13'd66,  13'd306,  -13'd5,  -13'd210,  13'd254,  13'd92,  -13'd360,  13'd201,  -13'd174,  13'd460,  13'd52,  -13'd173,  -13'd661,  -13'd521,  -13'd506,  13'd395,  
-13'd168,  13'd172,  13'd124,  13'd186,  -13'd1037,  13'd225,  -13'd19,  13'd53,  13'd1068,  13'd223,  13'd214,  13'd197,  -13'd519,  13'd260,  13'd524,  -13'd149,  
13'd135,  -13'd545,  13'd10,  13'd431,  13'd282,  -13'd429,  -13'd74,  13'd421,  13'd409,  13'd312,  13'd574,  13'd289,  -13'd74,  13'd180,  -13'd58,  -13'd140,  
13'd624,  -13'd696,  -13'd508,  13'd305,  -13'd34,  13'd653,  13'd630,  13'd612,  13'd240,  13'd285,  -13'd359,  13'd86,  13'd455,  -13'd820,  13'd482,  13'd685,  
13'd50,  13'd728,  13'd207,  -13'd534,  13'd428,  -13'd186,  13'd113,  13'd25,  -13'd6,  13'd354,  13'd31,  -13'd194,  -13'd374,  13'd329,  -13'd291,  -13'd159,  
13'd539,  -13'd526,  13'd568,  13'd99,  -13'd783,  13'd475,  -13'd117,  13'd259,  13'd521,  13'd1219,  -13'd276,  13'd293,  -13'd235,  13'd20,  -13'd443,  13'd581,  

13'd475,  -13'd707,  -13'd396,  -13'd244,  -13'd749,  13'd250,  13'd960,  -13'd709,  13'd498,  -13'd218,  -13'd98,  13'd570,  -13'd258,  -13'd45,  -13'd779,  -13'd808,  
-13'd470,  -13'd416,  -13'd949,  -13'd58,  -13'd1,  13'd322,  -13'd123,  -13'd341,  -13'd262,  13'd474,  -13'd437,  -13'd187,  -13'd579,  -13'd126,  13'd201,  -13'd68,  
-13'd556,  13'd121,  -13'd671,  -13'd305,  13'd908,  -13'd286,  -13'd885,  -13'd118,  -13'd64,  13'd141,  -13'd8,  -13'd339,  -13'd44,  -13'd1774,  -13'd112,  13'd408,  
-13'd511,  -13'd415,  -13'd582,  -13'd32,  13'd283,  -13'd67,  -13'd741,  13'd326,  13'd324,  13'd411,  -13'd727,  13'd207,  -13'd388,  -13'd198,  -13'd431,  13'd185,  
-13'd742,  -13'd614,  13'd494,  13'd49,  -13'd33,  -13'd78,  -13'd394,  -13'd281,  -13'd140,  13'd461,  -13'd547,  -13'd292,  13'd705,  -13'd15,  13'd326,  13'd163,  
13'd18,  13'd241,  -13'd194,  -13'd240,  -13'd1109,  13'd139,  13'd104,  13'd428,  13'd187,  13'd204,  13'd698,  -13'd46,  -13'd4,  -13'd231,  -13'd123,  13'd456,  
13'd364,  13'd345,  -13'd355,  -13'd329,  -13'd508,  13'd106,  13'd312,  -13'd200,  -13'd95,  13'd261,  -13'd532,  13'd289,  -13'd479,  13'd478,  13'd206,  13'd657,  
13'd459,  -13'd512,  -13'd821,  -13'd69,  13'd141,  13'd332,  13'd98,  -13'd87,  -13'd70,  13'd51,  -13'd378,  13'd70,  13'd640,  -13'd1038,  13'd516,  -13'd77,  
-13'd10,  -13'd465,  -13'd826,  -13'd45,  13'd150,  -13'd444,  13'd342,  -13'd129,  13'd210,  -13'd430,  13'd232,  13'd55,  13'd312,  -13'd102,  -13'd146,  13'd324,  
-13'd872,  13'd122,  13'd758,  13'd40,  13'd44,  -13'd162,  13'd7,  13'd143,  -13'd551,  -13'd260,  13'd505,  -13'd530,  13'd220,  -13'd161,  13'd224,  -13'd234,  
-13'd245,  -13'd31,  13'd402,  13'd184,  13'd243,  -13'd129,  -13'd923,  13'd986,  13'd480,  -13'd145,  -13'd1804,  -13'd447,  13'd452,  13'd703,  13'd607,  -13'd200,  
13'd113,  13'd330,  -13'd373,  13'd794,  13'd456,  13'd79,  -13'd544,  13'd332,  -13'd673,  -13'd345,  13'd419,  -13'd522,  13'd524,  13'd41,  13'd566,  -13'd295,  
13'd234,  13'd663,  -13'd869,  -13'd634,  13'd52,  13'd415,  13'd601,  -13'd296,  -13'd258,  -13'd329,  -13'd319,  13'd395,  -13'd63,  -13'd1137,  -13'd442,  -13'd53,  
-13'd405,  13'd332,  13'd245,  -13'd1188,  13'd465,  13'd199,  -13'd352,  13'd68,  -13'd158,  -13'd609,  -13'd91,  13'd153,  13'd16,  -13'd122,  -13'd509,  13'd645,  
13'd340,  13'd3,  13'd48,  -13'd500,  -13'd444,  13'd624,  -13'd212,  -13'd275,  13'd553,  13'd473,  13'd490,  -13'd137,  -13'd721,  13'd254,  -13'd9,  13'd351,  
-13'd64,  -13'd880,  -13'd270,  13'd873,  13'd654,  13'd514,  -13'd1084,  13'd91,  -13'd234,  -13'd46,  -13'd342,  13'd33,  13'd487,  13'd123,  13'd3,  -13'd251,  
-13'd152,  -13'd308,  -13'd52,  -13'd60,  13'd1138,  13'd153,  -13'd120,  -13'd244,  13'd60,  -13'd624,  13'd465,  -13'd131,  13'd574,  -13'd57,  -13'd85,  13'd6,  
13'd566,  13'd946,  13'd158,  -13'd96,  13'd913,  -13'd565,  13'd39,  13'd71,  -13'd672,  -13'd52,  13'd798,  -13'd477,  -13'd503,  13'd161,  -13'd474,  -13'd259,  
13'd320,  13'd552,  -13'd741,  -13'd277,  13'd788,  13'd621,  -13'd215,  -13'd213,  13'd636,  -13'd192,  -13'd509,  13'd658,  -13'd152,  13'd160,  -13'd472,  -13'd720,  
-13'd659,  -13'd1030,  13'd199,  -13'd413,  -13'd650,  13'd109,  -13'd116,  13'd131,  13'd724,  -13'd6,  -13'd290,  -13'd738,  13'd514,  13'd348,  -13'd172,  -13'd704,  
13'd5,  13'd469,  -13'd168,  13'd635,  13'd852,  13'd384,  -13'd98,  13'd16,  13'd264,  13'd658,  13'd86,  13'd494,  13'd199,  -13'd738,  13'd898,  13'd89,  
13'd75,  -13'd253,  13'd198,  13'd527,  13'd491,  -13'd741,  13'd178,  -13'd83,  13'd514,  -13'd697,  13'd339,  13'd60,  13'd137,  -13'd448,  13'd24,  -13'd351,  
13'd619,  13'd37,  13'd400,  13'd514,  13'd85,  13'd613,  -13'd119,  -13'd254,  13'd869,  13'd315,  13'd474,  13'd600,  -13'd7,  -13'd613,  -13'd341,  13'd161,  
13'd502,  13'd324,  -13'd45,  -13'd214,  13'd157,  -13'd207,  -13'd227,  -13'd319,  13'd694,  -13'd252,  -13'd431,  13'd384,  13'd599,  13'd97,  13'd385,  -13'd332,  
13'd1032,  -13'd519,  13'd741,  13'd273,  -13'd484,  13'd399,  13'd896,  -13'd293,  13'd1435,  13'd322,  -13'd130,  13'd1055,  13'd106,  13'd347,  13'd164,  -13'd422,  

-13'd442,  13'd418,  13'd556,  -13'd306,  13'd224,  13'd82,  13'd230,  13'd738,  13'd326,  -13'd263,  -13'd281,  13'd35,  13'd79,  13'd473,  -13'd541,  13'd967,  
-13'd137,  13'd526,  13'd951,  -13'd1125,  13'd136,  -13'd462,  13'd741,  13'd231,  -13'd381,  -13'd32,  13'd4,  13'd305,  13'd150,  13'd517,  13'd65,  -13'd303,  
-13'd422,  13'd51,  13'd248,  -13'd370,  13'd474,  -13'd794,  13'd396,  -13'd446,  -13'd70,  -13'd292,  13'd595,  13'd800,  13'd682,  13'd1541,  -13'd445,  13'd413,  
-13'd241,  13'd762,  13'd202,  -13'd321,  13'd639,  -13'd9,  13'd860,  13'd382,  -13'd57,  -13'd1095,  -13'd242,  -13'd45,  13'd241,  13'd1718,  -13'd311,  -13'd122,  
13'd474,  13'd205,  -13'd388,  -13'd141,  -13'd925,  13'd49,  13'd346,  -13'd284,  -13'd270,  -13'd327,  13'd115,  13'd252,  13'd568,  -13'd11,  -13'd284,  -13'd502,  
-13'd413,  -13'd130,  -13'd226,  13'd97,  13'd521,  -13'd420,  13'd52,  -13'd378,  -13'd533,  13'd439,  -13'd105,  -13'd484,  13'd70,  13'd768,  13'd287,  -13'd216,  
13'd604,  -13'd676,  13'd284,  13'd867,  -13'd298,  -13'd1,  13'd442,  -13'd24,  -13'd70,  -13'd380,  13'd535,  13'd253,  -13'd341,  13'd289,  -13'd475,  -13'd457,  
13'd731,  -13'd595,  13'd17,  13'd888,  -13'd36,  -13'd317,  13'd1037,  -13'd388,  -13'd715,  -13'd60,  -13'd133,  13'd172,  -13'd286,  -13'd655,  -13'd679,  -13'd1187,  
13'd1011,  13'd709,  13'd651,  -13'd329,  -13'd16,  13'd138,  -13'd76,  -13'd59,  13'd665,  13'd456,  -13'd255,  13'd176,  13'd217,  13'd292,  -13'd251,  -13'd582,  
13'd1155,  -13'd297,  -13'd320,  -13'd215,  13'd229,  -13'd77,  13'd504,  -13'd45,  13'd230,  13'd575,  -13'd79,  13'd526,  -13'd295,  -13'd94,  13'd73,  13'd182,  
-13'd350,  13'd98,  13'd451,  -13'd248,  13'd143,  13'd75,  13'd364,  13'd231,  -13'd39,  13'd128,  13'd305,  -13'd528,  -13'd300,  -13'd575,  -13'd436,  13'd770,  
13'd396,  13'd481,  -13'd130,  13'd711,  -13'd143,  -13'd315,  -13'd304,  13'd72,  -13'd335,  13'd325,  13'd312,  13'd208,  -13'd31,  13'd295,  13'd148,  -13'd120,  
-13'd72,  -13'd757,  -13'd351,  13'd109,  -13'd90,  13'd440,  -13'd380,  -13'd147,  -13'd110,  13'd110,  13'd140,  -13'd105,  -13'd49,  -13'd790,  -13'd175,  13'd504,  
-13'd190,  -13'd112,  13'd67,  13'd497,  13'd202,  13'd160,  -13'd11,  -13'd641,  13'd337,  13'd58,  -13'd0,  13'd636,  13'd58,  -13'd263,  -13'd36,  13'd795,  
-13'd362,  -13'd572,  13'd162,  13'd61,  13'd111,  13'd362,  -13'd286,  -13'd326,  13'd267,  13'd230,  13'd270,  13'd410,  -13'd162,  -13'd856,  13'd970,  13'd312,  
13'd229,  13'd602,  -13'd247,  -13'd238,  -13'd784,  -13'd181,  -13'd92,  -13'd61,  -13'd262,  -13'd167,  13'd396,  -13'd215,  13'd634,  -13'd51,  -13'd41,  13'd299,  
13'd60,  -13'd296,  13'd136,  13'd291,  13'd189,  13'd210,  -13'd197,  -13'd84,  -13'd125,  -13'd346,  -13'd846,  13'd500,  -13'd44,  -13'd236,  13'd237,  13'd84,  
13'd48,  13'd431,  -13'd246,  -13'd101,  13'd699,  13'd92,  -13'd345,  13'd533,  13'd125,  -13'd294,  13'd225,  13'd213,  -13'd417,  -13'd73,  -13'd371,  -13'd468,  
-13'd14,  -13'd191,  -13'd187,  13'd419,  -13'd213,  13'd285,  13'd597,  13'd97,  13'd121,  13'd2,  13'd327,  -13'd42,  13'd389,  -13'd332,  -13'd200,  13'd184,  
-13'd305,  13'd1158,  -13'd50,  13'd277,  13'd458,  -13'd170,  13'd188,  -13'd15,  -13'd414,  -13'd571,  13'd196,  -13'd100,  -13'd42,  13'd650,  -13'd569,  13'd58,  
-13'd113,  13'd244,  13'd327,  -13'd1134,  -13'd1184,  13'd137,  13'd516,  -13'd332,  13'd315,  13'd185,  -13'd484,  -13'd513,  13'd101,  13'd813,  -13'd529,  -13'd284,  
-13'd250,  13'd334,  13'd395,  -13'd349,  -13'd37,  13'd481,  13'd436,  13'd56,  13'd20,  13'd394,  -13'd442,  13'd821,  -13'd235,  13'd647,  -13'd206,  13'd121,  
-13'd304,  13'd436,  13'd41,  -13'd374,  -13'd177,  13'd494,  13'd171,  13'd294,  13'd119,  -13'd643,  -13'd37,  -13'd79,  13'd350,  13'd81,  -13'd42,  -13'd857,  
-13'd221,  -13'd64,  -13'd629,  -13'd127,  13'd115,  -13'd229,  13'd421,  -13'd518,  13'd40,  -13'd95,  13'd31,  -13'd393,  -13'd66,  13'd432,  -13'd89,  13'd368,  
13'd812,  -13'd554,  -13'd613,  -13'd755,  -13'd677,  -13'd136,  13'd169,  -13'd177,  -13'd566,  -13'd1192,  -13'd410,  -13'd1339,  -13'd132,  -13'd190,  -13'd393,  -13'd825,  

-13'd72,  -13'd379,  13'd147,  13'd125,  -13'd217,  -13'd289,  13'd1170,  -13'd379,  -13'd4,  -13'd45,  -13'd868,  13'd157,  -13'd1113,  -13'd497,  13'd106,  -13'd14,  
-13'd843,  -13'd331,  13'd123,  -13'd552,  -13'd230,  -13'd223,  -13'd163,  -13'd957,  -13'd841,  -13'd148,  13'd507,  -13'd657,  -13'd322,  13'd29,  -13'd34,  -13'd308,  
-13'd262,  -13'd288,  13'd127,  -13'd622,  13'd151,  -13'd446,  13'd198,  13'd291,  13'd268,  13'd150,  13'd435,  -13'd255,  13'd179,  -13'd706,  13'd233,  13'd102,  
-13'd199,  13'd309,  13'd249,  13'd907,  -13'd253,  13'd570,  -13'd111,  13'd583,  13'd491,  -13'd60,  -13'd139,  13'd100,  -13'd181,  13'd129,  -13'd116,  -13'd434,  
13'd217,  13'd167,  -13'd157,  13'd1082,  -13'd737,  13'd134,  -13'd394,  13'd160,  -13'd231,  -13'd21,  13'd105,  -13'd79,  13'd941,  13'd2,  13'd368,  -13'd101,  
-13'd127,  -13'd335,  -13'd255,  13'd350,  -13'd668,  -13'd332,  13'd567,  -13'd251,  13'd41,  13'd117,  13'd329,  -13'd603,  13'd80,  -13'd315,  13'd117,  -13'd47,  
13'd812,  -13'd578,  -13'd294,  13'd251,  -13'd326,  -13'd655,  -13'd50,  13'd245,  13'd488,  13'd94,  -13'd263,  -13'd35,  -13'd608,  13'd348,  13'd71,  -13'd674,  
-13'd34,  -13'd966,  -13'd244,  13'd156,  13'd585,  13'd85,  13'd86,  13'd157,  13'd908,  13'd603,  13'd528,  -13'd346,  13'd177,  -13'd8,  13'd765,  -13'd304,  
-13'd599,  13'd183,  -13'd266,  -13'd367,  13'd432,  -13'd547,  13'd75,  13'd893,  13'd364,  13'd16,  13'd321,  -13'd709,  13'd40,  -13'd1016,  13'd76,  13'd433,  
-13'd948,  -13'd922,  13'd292,  -13'd197,  13'd386,  13'd45,  -13'd1016,  13'd187,  13'd364,  13'd376,  -13'd0,  13'd35,  13'd792,  13'd189,  -13'd724,  -13'd30,  
-13'd143,  13'd228,  -13'd392,  13'd628,  13'd24,  13'd521,  -13'd47,  13'd573,  13'd165,  -13'd204,  -13'd1271,  -13'd433,  13'd33,  13'd723,  13'd390,  13'd108,  
13'd12,  13'd131,  13'd281,  -13'd39,  -13'd675,  -13'd289,  -13'd480,  13'd455,  -13'd307,  13'd135,  -13'd162,  -13'd536,  -13'd331,  13'd335,  13'd200,  -13'd549,  
-13'd718,  -13'd48,  -13'd651,  -13'd11,  13'd352,  13'd308,  -13'd159,  -13'd157,  -13'd432,  13'd103,  13'd194,  -13'd805,  13'd267,  13'd18,  -13'd586,  13'd601,  
-13'd1011,  -13'd359,  -13'd113,  -13'd317,  13'd441,  13'd520,  -13'd464,  13'd28,  13'd279,  13'd43,  13'd177,  -13'd481,  -13'd22,  -13'd686,  -13'd299,  13'd688,  
-13'd1237,  -13'd281,  13'd763,  13'd436,  13'd379,  -13'd746,  13'd510,  -13'd558,  -13'd380,  13'd448,  -13'd459,  13'd302,  -13'd806,  13'd105,  13'd378,  -13'd134,  
-13'd225,  13'd357,  13'd132,  13'd855,  13'd191,  13'd706,  -13'd220,  -13'd6,  -13'd58,  13'd321,  -13'd57,  -13'd739,  13'd378,  13'd733,  -13'd156,  13'd452,  
-13'd397,  13'd436,  -13'd75,  13'd235,  13'd1,  13'd411,  -13'd392,  -13'd248,  -13'd444,  -13'd403,  13'd588,  -13'd54,  -13'd119,  13'd120,  13'd96,  -13'd78,  
13'd400,  13'd11,  -13'd395,  13'd134,  -13'd402,  -13'd575,  13'd363,  13'd499,  -13'd577,  13'd363,  13'd591,  13'd266,  13'd244,  13'd24,  -13'd229,  -13'd277,  
13'd162,  13'd899,  -13'd6,  -13'd871,  13'd75,  13'd317,  13'd290,  13'd350,  13'd619,  -13'd1154,  -13'd20,  13'd446,  -13'd6,  13'd277,  -13'd307,  13'd238,  
13'd104,  13'd97,  13'd517,  -13'd479,  13'd313,  -13'd291,  13'd1040,  13'd1138,  -13'd38,  -13'd1127,  -13'd404,  13'd39,  13'd159,  13'd294,  13'd250,  -13'd663,  
13'd336,  13'd370,  -13'd804,  13'd296,  13'd1000,  13'd122,  13'd73,  13'd121,  13'd1211,  13'd467,  13'd224,  13'd377,  -13'd485,  -13'd962,  -13'd407,  13'd418,  
-13'd87,  13'd210,  -13'd950,  13'd698,  -13'd26,  13'd421,  13'd141,  -13'd132,  13'd504,  13'd594,  13'd689,  13'd98,  -13'd360,  -13'd672,  -13'd347,  13'd196,  
13'd779,  13'd438,  13'd368,  13'd441,  13'd348,  -13'd224,  13'd168,  -13'd390,  13'd976,  -13'd94,  13'd276,  13'd607,  13'd199,  13'd380,  -13'd33,  13'd193,  
13'd517,  13'd13,  13'd392,  -13'd810,  -13'd113,  -13'd349,  13'd247,  13'd382,  13'd178,  13'd668,  -13'd51,  13'd857,  13'd425,  13'd900,  13'd181,  -13'd176,  
13'd540,  13'd32,  -13'd404,  -13'd554,  -13'd644,  13'd505,  13'd185,  -13'd358,  -13'd103,  -13'd372,  -13'd175,  13'd295,  13'd422,  13'd779,  -13'd90,  -13'd221,  

-13'd1222,  13'd545,  13'd66,  -13'd726,  -13'd14,  13'd62,  13'd273,  -13'd848,  -13'd227,  -13'd856,  -13'd1068,  13'd192,  -13'd970,  13'd325,  -13'd498,  13'd424,  
-13'd412,  13'd132,  13'd862,  13'd38,  13'd408,  -13'd493,  -13'd213,  -13'd482,  -13'd419,  -13'd482,  -13'd593,  13'd380,  -13'd357,  13'd62,  -13'd471,  -13'd82,  
13'd178,  13'd1071,  -13'd161,  -13'd437,  13'd482,  13'd526,  -13'd528,  -13'd848,  13'd511,  13'd47,  -13'd179,  13'd259,  -13'd911,  13'd927,  -13'd76,  13'd217,  
13'd328,  13'd442,  -13'd305,  13'd63,  -13'd137,  13'd612,  -13'd29,  -13'd485,  13'd416,  -13'd151,  -13'd189,  -13'd383,  -13'd109,  13'd642,  -13'd330,  13'd400,  
13'd725,  13'd866,  -13'd929,  -13'd194,  13'd99,  13'd612,  13'd210,  -13'd294,  13'd57,  -13'd666,  13'd358,  13'd378,  13'd368,  -13'd320,  -13'd93,  -13'd152,  
13'd128,  13'd134,  13'd508,  -13'd116,  -13'd97,  -13'd22,  13'd402,  -13'd683,  -13'd1160,  13'd315,  -13'd187,  13'd831,  -13'd658,  13'd446,  13'd574,  -13'd588,  
13'd110,  -13'd618,  13'd231,  -13'd250,  13'd350,  -13'd332,  13'd140,  -13'd21,  13'd513,  13'd3,  -13'd220,  13'd853,  -13'd288,  13'd275,  -13'd124,  -13'd647,  
13'd183,  13'd164,  13'd281,  -13'd275,  13'd390,  -13'd459,  13'd384,  -13'd465,  -13'd398,  13'd181,  -13'd241,  -13'd583,  13'd735,  -13'd275,  13'd689,  -13'd847,  
-13'd141,  -13'd813,  13'd289,  -13'd256,  13'd799,  -13'd200,  13'd120,  13'd324,  -13'd242,  -13'd367,  -13'd1069,  13'd585,  -13'd747,  13'd38,  -13'd570,  13'd202,  
13'd263,  13'd529,  -13'd413,  -13'd608,  -13'd547,  -13'd249,  13'd461,  -13'd378,  13'd382,  -13'd279,  13'd711,  -13'd713,  -13'd68,  -13'd299,  -13'd59,  -13'd358,  
13'd102,  -13'd361,  13'd220,  13'd423,  -13'd751,  13'd84,  13'd118,  13'd278,  13'd287,  13'd444,  -13'd0,  -13'd245,  -13'd378,  13'd955,  13'd555,  -13'd450,  
-13'd21,  -13'd127,  13'd270,  13'd593,  -13'd403,  13'd771,  13'd161,  -13'd312,  13'd71,  13'd223,  -13'd600,  13'd296,  13'd505,  -13'd379,  -13'd129,  13'd268,  
13'd339,  -13'd191,  -13'd493,  13'd893,  13'd64,  -13'd90,  -13'd190,  13'd385,  -13'd580,  -13'd382,  13'd516,  -13'd471,  13'd492,  13'd294,  13'd714,  13'd441,  
13'd494,  -13'd326,  13'd1035,  13'd199,  -13'd526,  13'd897,  13'd427,  13'd309,  13'd67,  -13'd660,  13'd47,  13'd132,  -13'd25,  -13'd263,  13'd116,  -13'd92,  
-13'd271,  -13'd284,  -13'd545,  13'd33,  -13'd75,  13'd129,  13'd66,  13'd141,  -13'd589,  -13'd343,  13'd155,  -13'd247,  13'd617,  13'd406,  -13'd176,  13'd318,  
13'd576,  -13'd419,  -13'd277,  13'd406,  13'd508,  13'd129,  13'd197,  13'd47,  -13'd597,  13'd311,  13'd431,  -13'd10,  13'd267,  13'd594,  13'd439,  13'd563,  
-13'd855,  13'd395,  13'd60,  13'd86,  13'd705,  -13'd542,  13'd385,  -13'd179,  13'd190,  13'd6,  13'd314,  13'd211,  13'd228,  -13'd157,  -13'd568,  13'd370,  
-13'd132,  13'd48,  -13'd249,  13'd342,  13'd14,  -13'd359,  -13'd112,  13'd138,  -13'd203,  -13'd22,  -13'd429,  -13'd585,  -13'd75,  -13'd449,  13'd357,  -13'd100,  
-13'd384,  13'd22,  -13'd315,  -13'd124,  -13'd22,  -13'd136,  -13'd189,  13'd835,  -13'd876,  -13'd369,  13'd286,  13'd291,  -13'd424,  -13'd666,  -13'd186,  -13'd375,  
13'd356,  -13'd442,  -13'd1215,  -13'd17,  -13'd767,  13'd341,  -13'd263,  13'd181,  -13'd407,  -13'd423,  13'd102,  -13'd18,  -13'd168,  -13'd578,  13'd347,  13'd588,  
-13'd83,  13'd610,  13'd628,  13'd69,  13'd580,  13'd452,  -13'd137,  13'd573,  -13'd336,  -13'd549,  13'd330,  13'd478,  -13'd122,  -13'd423,  13'd50,  13'd38,  
13'd392,  13'd146,  13'd369,  -13'd162,  13'd665,  -13'd278,  13'd138,  -13'd471,  -13'd40,  -13'd105,  -13'd145,  -13'd178,  13'd4,  13'd313,  -13'd712,  13'd251,  
-13'd238,  13'd146,  -13'd377,  -13'd729,  13'd142,  -13'd630,  -13'd117,  -13'd301,  -13'd560,  13'd664,  -13'd258,  -13'd145,  -13'd122,  13'd672,  13'd202,  -13'd240,  
-13'd246,  13'd168,  13'd551,  13'd538,  13'd664,  -13'd521,  -13'd99,  -13'd111,  -13'd155,  13'd257,  13'd106,  13'd489,  13'd13,  13'd129,  -13'd234,  -13'd66,  
-13'd387,  -13'd569,  13'd239,  13'd844,  13'd227,  13'd213,  13'd317,  -13'd332,  -13'd581,  13'd796,  -13'd207,  13'd235,  -13'd256,  -13'd792,  13'd49,  13'd166,  

13'd8,  -13'd534,  -13'd145,  13'd301,  -13'd138,  -13'd79,  13'd80,  13'd284,  -13'd166,  -13'd83,  13'd1209,  -13'd596,  13'd498,  -13'd282,  13'd139,  13'd726,  
13'd408,  -13'd26,  13'd201,  -13'd81,  -13'd346,  13'd645,  13'd89,  13'd97,  13'd35,  -13'd575,  13'd1056,  -13'd21,  -13'd464,  -13'd622,  -13'd715,  -13'd336,  
-13'd189,  13'd327,  13'd375,  13'd210,  -13'd149,  -13'd295,  -13'd190,  -13'd330,  -13'd558,  -13'd612,  13'd608,  13'd277,  -13'd71,  -13'd115,  13'd6,  13'd791,  
13'd1008,  -13'd189,  -13'd774,  -13'd192,  -13'd185,  -13'd423,  -13'd512,  13'd548,  13'd356,  13'd550,  13'd515,  -13'd104,  13'd19,  -13'd802,  -13'd40,  13'd91,  
13'd77,  13'd127,  13'd489,  13'd739,  -13'd165,  13'd409,  -13'd71,  13'd413,  13'd589,  13'd426,  13'd21,  -13'd139,  -13'd285,  13'd235,  13'd306,  13'd23,  
-13'd812,  13'd360,  13'd814,  13'd259,  13'd3,  -13'd596,  13'd89,  -13'd238,  -13'd286,  13'd273,  -13'd225,  13'd391,  -13'd1055,  -13'd599,  13'd615,  13'd522,  
-13'd463,  13'd211,  -13'd281,  -13'd420,  -13'd167,  -13'd144,  13'd830,  -13'd568,  13'd247,  -13'd159,  13'd915,  -13'd134,  13'd145,  -13'd276,  -13'd1073,  -13'd70,  
-13'd253,  13'd999,  13'd38,  13'd41,  13'd104,  13'd265,  13'd720,  -13'd599,  -13'd261,  -13'd116,  13'd395,  -13'd394,  13'd169,  13'd648,  -13'd1025,  13'd1,  
-13'd365,  13'd488,  -13'd320,  -13'd259,  13'd523,  13'd283,  -13'd517,  13'd53,  13'd457,  -13'd43,  13'd798,  -13'd481,  13'd402,  13'd475,  13'd470,  13'd220,  
-13'd617,  -13'd669,  -13'd614,  13'd134,  13'd302,  -13'd202,  13'd309,  -13'd494,  13'd109,  -13'd129,  -13'd479,  -13'd141,  -13'd249,  13'd92,  13'd776,  -13'd59,  
13'd202,  -13'd428,  13'd318,  -13'd469,  -13'd592,  13'd623,  13'd91,  13'd304,  13'd201,  -13'd316,  -13'd871,  13'd218,  13'd4,  -13'd425,  13'd305,  -13'd235,  
13'd639,  -13'd40,  -13'd108,  13'd398,  13'd550,  13'd612,  -13'd292,  -13'd135,  13'd435,  13'd149,  13'd106,  -13'd105,  13'd81,  -13'd449,  13'd50,  -13'd21,  
13'd415,  -13'd178,  13'd65,  -13'd691,  -13'd291,  -13'd100,  -13'd438,  -13'd118,  13'd155,  13'd812,  -13'd406,  -13'd462,  13'd524,  13'd227,  -13'd756,  -13'd223,  
13'd564,  -13'd379,  -13'd44,  -13'd77,  13'd518,  13'd670,  13'd140,  -13'd525,  -13'd139,  -13'd512,  -13'd66,  13'd265,  -13'd1549,  13'd590,  -13'd292,  13'd57,  
13'd194,  13'd264,  13'd1318,  -13'd344,  -13'd808,  13'd41,  13'd818,  13'd352,  13'd507,  13'd602,  -13'd731,  13'd1139,  -13'd700,  -13'd182,  -13'd482,  -13'd28,  
13'd625,  13'd636,  13'd651,  -13'd508,  -13'd632,  -13'd3,  -13'd174,  13'd627,  -13'd72,  -13'd195,  -13'd743,  13'd110,  -13'd174,  -13'd38,  -13'd157,  13'd94,  
-13'd178,  -13'd42,  13'd669,  13'd275,  -13'd555,  -13'd666,  13'd739,  -13'd253,  13'd264,  -13'd50,  13'd614,  13'd628,  13'd297,  13'd153,  -13'd138,  -13'd182,  
-13'd763,  -13'd356,  13'd612,  -13'd17,  -13'd496,  -13'd145,  13'd104,  -13'd53,  -13'd124,  13'd325,  13'd266,  13'd109,  -13'd221,  13'd612,  -13'd80,  13'd39,  
13'd901,  13'd584,  -13'd195,  13'd14,  -13'd678,  -13'd667,  13'd527,  13'd14,  13'd302,  13'd342,  13'd268,  13'd628,  13'd681,  13'd121,  -13'd188,  13'd100,  
13'd428,  13'd181,  13'd303,  13'd247,  13'd359,  13'd314,  -13'd324,  13'd554,  13'd639,  -13'd457,  13'd352,  13'd800,  13'd111,  13'd451,  13'd407,  13'd604,  
-13'd491,  13'd345,  13'd130,  -13'd500,  -13'd1077,  13'd484,  13'd186,  13'd285,  -13'd1040,  -13'd15,  -13'd241,  13'd502,  -13'd626,  13'd693,  -13'd648,  13'd436,  
13'd389,  13'd657,  -13'd493,  -13'd363,  -13'd78,  -13'd470,  13'd392,  -13'd127,  13'd731,  -13'd341,  -13'd357,  13'd11,  13'd323,  13'd530,  13'd821,  13'd242,  
-13'd406,  13'd116,  13'd438,  -13'd754,  -13'd406,  13'd131,  13'd283,  13'd260,  -13'd514,  -13'd222,  -13'd177,  -13'd437,  13'd407,  -13'd358,  13'd79,  13'd318,  
13'd77,  -13'd302,  13'd858,  -13'd222,  -13'd499,  -13'd789,  13'd568,  -13'd340,  -13'd268,  -13'd293,  13'd203,  -13'd98,  -13'd600,  13'd512,  -13'd40,  -13'd387,  
-13'd760,  -13'd322,  -13'd923,  -13'd692,  13'd36,  -13'd75,  -13'd294,  13'd138,  -13'd1194,  -13'd586,  -13'd579,  -13'd1079,  -13'd382,  13'd336,  -13'd653,  -13'd114,  

13'd82,  13'd187,  -13'd180,  13'd21,  13'd237,  13'd71,  -13'd13,  13'd769,  13'd92,  -13'd575,  13'd601,  -13'd45,  -13'd238,  -13'd218,  -13'd551,  -13'd342,  
13'd178,  13'd287,  13'd10,  13'd132,  13'd85,  13'd275,  13'd415,  13'd15,  -13'd492,  -13'd975,  -13'd751,  13'd181,  -13'd98,  13'd774,  13'd449,  13'd114,  
13'd604,  13'd298,  -13'd316,  13'd258,  -13'd406,  13'd98,  -13'd192,  -13'd648,  13'd779,  -13'd804,  -13'd297,  13'd447,  -13'd188,  13'd447,  -13'd95,  13'd79,  
-13'd235,  13'd177,  13'd398,  -13'd877,  13'd221,  -13'd95,  -13'd1,  13'd247,  13'd21,  13'd797,  13'd113,  -13'd11,  13'd450,  13'd768,  -13'd753,  13'd747,  
13'd97,  13'd334,  13'd176,  13'd205,  13'd159,  13'd231,  13'd518,  -13'd456,  13'd369,  13'd241,  13'd496,  13'd342,  13'd345,  -13'd700,  -13'd170,  13'd39,  
13'd71,  -13'd309,  -13'd982,  13'd527,  -13'd91,  -13'd57,  13'd153,  -13'd767,  -13'd3,  -13'd88,  -13'd371,  13'd78,  -13'd360,  -13'd341,  -13'd733,  -13'd183,  
13'd262,  13'd169,  13'd802,  13'd17,  -13'd618,  -13'd351,  -13'd726,  -13'd20,  -13'd258,  13'd30,  13'd438,  13'd418,  -13'd581,  13'd195,  13'd181,  13'd359,  
-13'd589,  -13'd716,  13'd322,  13'd448,  13'd130,  -13'd163,  -13'd337,  -13'd218,  -13'd237,  -13'd228,  13'd159,  -13'd234,  -13'd861,  -13'd50,  13'd661,  -13'd148,  
-13'd604,  13'd361,  -13'd117,  -13'd202,  -13'd23,  -13'd133,  -13'd169,  13'd43,  13'd173,  -13'd277,  -13'd529,  13'd238,  -13'd147,  13'd235,  13'd223,  -13'd241,  
13'd180,  13'd915,  13'd80,  13'd47,  -13'd99,  -13'd405,  -13'd187,  -13'd402,  13'd158,  13'd618,  -13'd740,  13'd633,  13'd157,  -13'd247,  -13'd309,  13'd476,  
13'd479,  13'd782,  -13'd607,  13'd114,  -13'd773,  13'd471,  -13'd195,  -13'd454,  13'd347,  -13'd438,  13'd649,  -13'd21,  -13'd36,  13'd72,  13'd703,  -13'd564,  
13'd225,  13'd503,  -13'd157,  13'd213,  -13'd142,  -13'd72,  -13'd152,  -13'd203,  13'd782,  13'd713,  13'd25,  13'd627,  13'd962,  13'd382,  -13'd785,  13'd55,  
-13'd117,  -13'd182,  -13'd19,  -13'd363,  -13'd311,  -13'd207,  13'd110,  13'd46,  13'd723,  -13'd67,  13'd88,  13'd416,  13'd381,  13'd4,  -13'd529,  -13'd271,  
-13'd338,  -13'd405,  13'd223,  13'd323,  -13'd421,  -13'd193,  -13'd344,  13'd60,  -13'd227,  13'd304,  -13'd547,  13'd272,  13'd304,  13'd558,  13'd69,  -13'd423,  
13'd872,  -13'd101,  -13'd965,  13'd220,  13'd162,  13'd951,  -13'd702,  -13'd131,  13'd658,  -13'd219,  13'd293,  -13'd122,  13'd236,  13'd330,  -13'd284,  13'd166,  
13'd769,  -13'd127,  13'd847,  13'd304,  -13'd384,  -13'd330,  13'd118,  -13'd307,  13'd82,  -13'd388,  -13'd417,  13'd52,  13'd416,  13'd479,  -13'd232,  13'd85,  
13'd813,  13'd541,  -13'd75,  13'd4,  -13'd294,  -13'd789,  -13'd33,  13'd55,  13'd538,  13'd92,  13'd113,  13'd846,  13'd619,  13'd237,  -13'd99,  13'd3,  
-13'd93,  13'd154,  -13'd275,  13'd95,  13'd218,  13'd462,  13'd121,  13'd337,  13'd430,  -13'd708,  13'd231,  -13'd254,  13'd434,  -13'd415,  -13'd428,  13'd287,  
-13'd204,  -13'd57,  -13'd53,  13'd716,  13'd1047,  13'd495,  13'd299,  13'd192,  -13'd763,  13'd232,  -13'd162,  -13'd69,  -13'd518,  -13'd393,  13'd942,  13'd227,  
-13'd159,  -13'd482,  -13'd410,  13'd225,  -13'd425,  13'd132,  -13'd364,  13'd142,  -13'd177,  13'd1048,  13'd712,  13'd657,  13'd456,  13'd568,  -13'd70,  13'd372,  
-13'd1,  -13'd496,  13'd715,  13'd185,  -13'd3,  13'd187,  13'd365,  13'd469,  -13'd373,  13'd69,  -13'd245,  -13'd772,  13'd28,  13'd733,  13'd630,  13'd64,  
-13'd236,  -13'd98,  -13'd508,  -13'd172,  -13'd105,  13'd133,  13'd456,  13'd253,  -13'd301,  -13'd714,  13'd86,  13'd236,  -13'd47,  -13'd310,  -13'd328,  -13'd351,  
-13'd492,  -13'd180,  13'd39,  13'd289,  13'd357,  -13'd327,  -13'd702,  -13'd25,  -13'd1169,  -13'd536,  13'd454,  -13'd104,  -13'd371,  -13'd297,  -13'd436,  13'd148,  
-13'd967,  13'd117,  -13'd185,  13'd4,  -13'd14,  -13'd150,  -13'd191,  13'd261,  -13'd700,  13'd201,  -13'd372,  13'd104,  -13'd18,  -13'd391,  13'd64,  -13'd297,  
-13'd679,  -13'd101,  -13'd696,  13'd473,  13'd152,  -13'd239,  -13'd264,  13'd407,  13'd376,  13'd650,  13'd936,  13'd589,  13'd84,  13'd96,  13'd8,  13'd907,  

13'd351,  13'd436,  -13'd247,  -13'd459,  -13'd317,  -13'd244,  13'd105,  -13'd582,  -13'd480,  13'd1,  -13'd14,  13'd41,  -13'd529,  -13'd877,  -13'd633,  -13'd165,  
13'd614,  13'd240,  -13'd603,  13'd420,  -13'd529,  13'd226,  -13'd575,  13'd206,  13'd377,  -13'd189,  13'd396,  -13'd658,  -13'd80,  13'd38,  -13'd11,  -13'd35,  
13'd692,  -13'd342,  -13'd1076,  13'd705,  -13'd364,  -13'd331,  -13'd293,  -13'd168,  13'd770,  13'd326,  -13'd606,  13'd213,  13'd336,  -13'd1177,  -13'd124,  13'd1026,  
-13'd218,  -13'd452,  13'd204,  -13'd212,  13'd633,  -13'd199,  -13'd871,  13'd92,  13'd12,  13'd648,  -13'd753,  -13'd107,  13'd123,  13'd225,  13'd385,  13'd386,  
-13'd57,  13'd25,  13'd498,  13'd167,  13'd476,  -13'd118,  -13'd837,  -13'd17,  -13'd380,  13'd479,  -13'd912,  -13'd217,  -13'd270,  13'd42,  -13'd454,  -13'd297,  
13'd230,  13'd56,  13'd259,  -13'd129,  13'd57,  13'd249,  -13'd304,  13'd126,  -13'd7,  13'd299,  -13'd231,  13'd489,  -13'd396,  13'd126,  -13'd286,  13'd210,  
-13'd146,  13'd515,  -13'd548,  -13'd227,  -13'd218,  -13'd344,  -13'd608,  13'd706,  -13'd228,  13'd278,  -13'd909,  13'd171,  13'd373,  13'd741,  13'd336,  13'd596,  
-13'd366,  -13'd612,  13'd281,  -13'd265,  13'd415,  13'd94,  -13'd358,  13'd205,  13'd73,  13'd500,  -13'd377,  13'd369,  -13'd111,  -13'd167,  13'd530,  -13'd273,  
-13'd140,  -13'd220,  13'd214,  13'd53,  -13'd509,  13'd193,  13'd156,  -13'd394,  -13'd580,  -13'd872,  -13'd251,  -13'd353,  13'd376,  13'd189,  13'd172,  -13'd256,  
13'd101,  -13'd228,  13'd77,  13'd540,  -13'd480,  -13'd159,  13'd177,  -13'd367,  13'd283,  -13'd1065,  -13'd455,  -13'd204,  13'd339,  13'd151,  13'd130,  13'd100,  
13'd361,  13'd119,  -13'd438,  13'd184,  13'd877,  13'd352,  -13'd328,  -13'd185,  13'd422,  13'd848,  -13'd98,  13'd333,  13'd545,  13'd86,  13'd159,  -13'd391,  
-13'd409,  13'd314,  13'd595,  13'd188,  13'd99,  13'd619,  -13'd446,  13'd993,  -13'd406,  13'd354,  13'd170,  -13'd32,  13'd528,  13'd87,  13'd183,  -13'd128,  
13'd156,  13'd237,  13'd651,  -13'd3,  13'd254,  13'd58,  13'd856,  13'd319,  -13'd93,  -13'd385,  13'd5,  -13'd14,  13'd65,  13'd36,  13'd735,  -13'd598,  
13'd932,  13'd78,  13'd819,  -13'd88,  -13'd240,  13'd672,  13'd1010,  -13'd235,  -13'd391,  -13'd48,  13'd538,  -13'd701,  -13'd394,  13'd607,  -13'd441,  -13'd116,  
13'd1156,  13'd288,  -13'd1013,  13'd170,  -13'd774,  13'd386,  13'd8,  13'd243,  -13'd100,  -13'd886,  -13'd638,  -13'd369,  13'd910,  13'd527,  -13'd138,  13'd606,  
-13'd836,  -13'd106,  -13'd670,  13'd198,  13'd1565,  13'd585,  -13'd739,  -13'd337,  13'd76,  -13'd87,  -13'd315,  13'd317,  -13'd130,  -13'd648,  13'd367,  -13'd207,  
-13'd568,  13'd331,  13'd419,  13'd275,  13'd733,  -13'd222,  13'd50,  -13'd1,  -13'd52,  13'd301,  13'd460,  13'd97,  -13'd173,  13'd288,  -13'd941,  13'd280,  
13'd685,  -13'd402,  13'd472,  13'd177,  13'd162,  13'd434,  -13'd35,  13'd364,  13'd387,  -13'd128,  -13'd399,  13'd387,  -13'd138,  13'd194,  -13'd970,  -13'd195,  
-13'd253,  13'd342,  13'd437,  -13'd490,  -13'd66,  -13'd574,  13'd496,  -13'd329,  -13'd113,  13'd439,  -13'd579,  -13'd123,  -13'd594,  13'd553,  -13'd69,  13'd401,  
-13'd229,  -13'd403,  13'd104,  13'd552,  -13'd345,  -13'd252,  -13'd565,  -13'd163,  13'd123,  -13'd121,  -13'd771,  -13'd688,  -13'd360,  13'd902,  -13'd205,  -13'd329,  
-13'd185,  13'd55,  -13'd333,  13'd349,  13'd714,  -13'd358,  -13'd142,  -13'd295,  13'd450,  -13'd185,  13'd41,  -13'd165,  13'd185,  13'd20,  13'd243,  13'd133,  
-13'd332,  -13'd646,  -13'd0,  13'd618,  13'd179,  -13'd142,  13'd790,  13'd619,  13'd875,  13'd284,  13'd685,  -13'd478,  13'd23,  13'd118,  13'd110,  13'd396,  
-13'd446,  13'd81,  13'd47,  13'd305,  -13'd113,  -13'd40,  -13'd308,  -13'd621,  -13'd249,  -13'd147,  13'd11,  13'd48,  13'd86,  13'd379,  -13'd318,  13'd441,  
-13'd429,  -13'd686,  13'd184,  -13'd203,  13'd248,  -13'd42,  13'd295,  13'd448,  13'd303,  13'd151,  -13'd23,  -13'd569,  13'd75,  13'd400,  13'd452,  13'd516,  
-13'd176,  -13'd771,  13'd251,  -13'd22,  -13'd373,  13'd343,  -13'd26,  -13'd751,  13'd226,  -13'd216,  -13'd323,  13'd645,  13'd649,  13'd681,  13'd451,  13'd111,  

-13'd47,  13'd9,  -13'd600,  -13'd102,  -13'd7,  -13'd115,  -13'd202,  -13'd48,  -13'd682,  13'd175,  13'd379,  -13'd396,  -13'd69,  13'd380,  -13'd410,  13'd52,  
13'd125,  13'd85,  -13'd375,  13'd558,  -13'd251,  -13'd285,  13'd280,  -13'd522,  13'd613,  -13'd481,  13'd458,  -13'd700,  13'd480,  13'd122,  13'd278,  -13'd148,  
-13'd242,  13'd152,  -13'd322,  -13'd506,  -13'd240,  13'd361,  -13'd718,  -13'd441,  -13'd515,  13'd616,  -13'd606,  -13'd315,  13'd108,  -13'd72,  -13'd0,  -13'd150,  
-13'd305,  -13'd280,  -13'd194,  -13'd224,  -13'd100,  -13'd221,  -13'd364,  -13'd194,  -13'd325,  13'd425,  13'd453,  -13'd328,  -13'd87,  -13'd4,  13'd33,  13'd268,  
13'd14,  -13'd542,  -13'd24,  13'd344,  13'd427,  13'd257,  -13'd237,  13'd320,  13'd389,  13'd176,  13'd521,  -13'd295,  13'd364,  -13'd480,  -13'd49,  13'd372,  
13'd243,  -13'd90,  -13'd47,  13'd371,  -13'd410,  -13'd652,  -13'd234,  -13'd281,  13'd304,  13'd730,  13'd201,  13'd244,  13'd25,  -13'd69,  13'd638,  -13'd172,  
-13'd176,  -13'd71,  -13'd300,  -13'd250,  -13'd49,  -13'd746,  -13'd45,  13'd226,  -13'd30,  13'd170,  -13'd126,  -13'd303,  13'd289,  -13'd177,  -13'd317,  -13'd289,  
-13'd418,  13'd667,  -13'd100,  13'd129,  13'd428,  13'd134,  13'd145,  13'd66,  -13'd381,  13'd30,  -13'd77,  -13'd369,  -13'd273,  -13'd376,  -13'd100,  -13'd407,  
13'd555,  -13'd48,  13'd557,  13'd203,  13'd213,  -13'd567,  -13'd436,  -13'd86,  13'd273,  -13'd408,  -13'd104,  -13'd558,  13'd192,  13'd483,  -13'd229,  -13'd591,  
13'd235,  13'd361,  13'd42,  13'd485,  -13'd32,  -13'd277,  -13'd525,  -13'd378,  -13'd731,  13'd181,  -13'd495,  -13'd345,  -13'd413,  13'd313,  -13'd167,  13'd372,  
13'd536,  -13'd854,  13'd338,  -13'd677,  -13'd236,  13'd415,  13'd163,  -13'd485,  -13'd265,  13'd184,  -13'd99,  -13'd359,  13'd443,  -13'd267,  -13'd244,  -13'd375,  
13'd714,  -13'd16,  -13'd129,  -13'd200,  -13'd202,  -13'd270,  13'd483,  -13'd103,  -13'd166,  -13'd249,  -13'd355,  -13'd51,  13'd171,  13'd212,  13'd284,  -13'd809,  
13'd523,  13'd290,  13'd103,  -13'd757,  13'd131,  13'd129,  -13'd843,  13'd70,  13'd70,  13'd595,  13'd395,  -13'd65,  13'd64,  13'd39,  13'd18,  13'd386,  
-13'd259,  13'd583,  -13'd667,  -13'd3,  -13'd430,  -13'd74,  -13'd312,  13'd271,  -13'd238,  13'd262,  13'd522,  -13'd518,  -13'd145,  -13'd200,  -13'd30,  13'd357,  
-13'd383,  -13'd71,  -13'd534,  -13'd800,  -13'd301,  13'd430,  -13'd188,  -13'd162,  13'd258,  -13'd72,  13'd229,  -13'd297,  -13'd193,  13'd94,  -13'd280,  -13'd585,  
-13'd307,  13'd108,  13'd92,  -13'd452,  13'd192,  -13'd508,  13'd665,  13'd335,  -13'd540,  13'd148,  13'd45,  13'd374,  -13'd148,  13'd19,  -13'd88,  -13'd244,  
13'd635,  13'd273,  13'd113,  -13'd454,  -13'd336,  -13'd215,  13'd408,  -13'd600,  13'd367,  -13'd17,  -13'd220,  -13'd326,  -13'd243,  -13'd575,  13'd71,  -13'd453,  
-13'd223,  -13'd173,  -13'd508,  13'd682,  -13'd62,  13'd751,  -13'd247,  -13'd371,  -13'd644,  13'd48,  -13'd634,  -13'd384,  -13'd369,  -13'd273,  -13'd356,  -13'd359,  
-13'd196,  13'd243,  13'd246,  13'd20,  -13'd125,  -13'd670,  13'd62,  13'd576,  13'd180,  -13'd317,  -13'd112,  13'd12,  13'd174,  -13'd136,  13'd180,  13'd387,  
-13'd534,  -13'd318,  13'd518,  13'd127,  -13'd14,  -13'd154,  -13'd294,  -13'd286,  -13'd643,  13'd309,  13'd267,  13'd354,  13'd620,  -13'd54,  -13'd452,  13'd208,  
-13'd119,  -13'd457,  13'd444,  13'd544,  -13'd190,  -13'd34,  -13'd846,  13'd498,  -13'd340,  -13'd368,  -13'd616,  -13'd418,  -13'd62,  -13'd408,  -13'd319,  -13'd385,  
-13'd21,  -13'd519,  -13'd46,  13'd8,  -13'd660,  -13'd156,  -13'd670,  -13'd91,  -13'd30,  -13'd271,  13'd622,  -13'd275,  -13'd653,  13'd95,  -13'd277,  -13'd285,  
-13'd604,  -13'd258,  13'd18,  13'd53,  13'd42,  -13'd454,  -13'd47,  -13'd626,  -13'd493,  13'd237,  -13'd430,  13'd483,  13'd35,  -13'd293,  13'd579,  -13'd537,  
13'd81,  13'd32,  -13'd114,  13'd501,  -13'd185,  13'd207,  -13'd309,  13'd306,  -13'd207,  -13'd295,  -13'd144,  -13'd365,  13'd218,  -13'd809,  -13'd67,  -13'd693,  
13'd537,  -13'd276,  -13'd450,  -13'd695,  -13'd255,  13'd392,  -13'd135,  -13'd53,  -13'd237,  -13'd215,  13'd137,  13'd194,  13'd488,  -13'd539,  13'd354,  13'd293,  

-13'd138,  13'd92,  13'd504,  13'd149,  -13'd409,  -13'd374,  13'd324,  13'd627,  13'd140,  13'd119,  -13'd8,  -13'd213,  13'd439,  13'd537,  -13'd2,  13'd188,  
-13'd288,  13'd89,  13'd1326,  -13'd997,  13'd569,  -13'd652,  13'd535,  13'd12,  -13'd365,  13'd66,  -13'd1304,  13'd158,  -13'd5,  13'd1031,  -13'd97,  13'd115,  
13'd232,  13'd157,  13'd0,  -13'd754,  13'd38,  -13'd484,  13'd1151,  13'd171,  -13'd350,  13'd11,  -13'd414,  -13'd171,  -13'd644,  13'd1354,  -13'd501,  -13'd735,  
-13'd443,  13'd381,  13'd366,  -13'd296,  13'd467,  -13'd236,  13'd709,  -13'd498,  13'd164,  -13'd180,  13'd119,  -13'd321,  -13'd751,  13'd701,  13'd548,  -13'd573,  
13'd582,  13'd507,  -13'd489,  -13'd187,  13'd16,  13'd1101,  13'd228,  13'd129,  13'd382,  13'd176,  13'd117,  -13'd255,  13'd243,  -13'd220,  -13'd129,  13'd224,  
13'd19,  -13'd232,  13'd36,  13'd297,  13'd270,  13'd90,  13'd220,  -13'd92,  -13'd618,  -13'd308,  -13'd360,  13'd443,  13'd79,  13'd364,  13'd81,  -13'd313,  
13'd639,  -13'd707,  13'd222,  13'd259,  -13'd272,  -13'd728,  13'd546,  -13'd21,  -13'd102,  -13'd341,  -13'd520,  13'd299,  -13'd702,  13'd1006,  -13'd594,  -13'd860,  
13'd39,  13'd511,  13'd588,  -13'd163,  -13'd473,  -13'd320,  13'd393,  -13'd305,  13'd300,  13'd41,  -13'd186,  -13'd98,  -13'd371,  13'd785,  13'd271,  -13'd957,  
13'd384,  -13'd94,  -13'd262,  -13'd827,  13'd551,  -13'd462,  -13'd179,  -13'd119,  -13'd227,  -13'd958,  -13'd235,  13'd256,  13'd240,  13'd348,  -13'd734,  -13'd63,  
13'd705,  13'd137,  13'd189,  -13'd478,  13'd52,  13'd572,  13'd170,  -13'd313,  13'd890,  13'd83,  13'd322,  -13'd226,  -13'd313,  -13'd110,  -13'd255,  -13'd325,  
-13'd359,  -13'd334,  -13'd907,  13'd205,  -13'd502,  13'd61,  13'd223,  -13'd400,  -13'd123,  -13'd313,  13'd995,  13'd222,  13'd714,  13'd317,  13'd219,  -13'd383,  
13'd182,  13'd71,  13'd65,  13'd137,  -13'd817,  13'd125,  13'd484,  -13'd493,  -13'd84,  13'd535,  -13'd218,  -13'd399,  13'd657,  13'd211,  13'd209,  13'd661,  
-13'd340,  13'd148,  13'd167,  13'd625,  13'd493,  13'd18,  13'd22,  -13'd72,  -13'd211,  -13'd308,  13'd537,  -13'd189,  13'd626,  -13'd321,  -13'd20,  -13'd190,  
-13'd319,  -13'd829,  13'd310,  13'd206,  13'd418,  13'd411,  13'd255,  13'd247,  13'd653,  -13'd469,  13'd42,  -13'd171,  -13'd272,  -13'd767,  -13'd74,  13'd277,  
-13'd429,  -13'd49,  -13'd530,  13'd505,  -13'd120,  13'd120,  -13'd66,  -13'd542,  -13'd660,  13'd505,  13'd106,  -13'd141,  13'd412,  -13'd516,  -13'd55,  13'd261,  
-13'd472,  13'd75,  13'd374,  -13'd553,  -13'd444,  -13'd295,  -13'd512,  -13'd19,  13'd362,  -13'd163,  13'd104,  13'd115,  13'd890,  -13'd18,  13'd421,  -13'd273,  
13'd117,  -13'd225,  -13'd41,  -13'd100,  13'd119,  13'd45,  13'd407,  13'd520,  -13'd302,  13'd215,  13'd686,  13'd672,  -13'd110,  13'd320,  -13'd287,  13'd165,  
13'd383,  -13'd628,  -13'd637,  13'd643,  13'd61,  13'd822,  -13'd182,  -13'd114,  -13'd658,  -13'd373,  13'd240,  13'd144,  13'd47,  13'd295,  13'd339,  -13'd81,  
-13'd16,  13'd50,  13'd412,  13'd702,  -13'd298,  13'd72,  13'd89,  13'd863,  13'd268,  13'd540,  13'd514,  13'd353,  -13'd366,  -13'd75,  13'd531,  13'd401,  
13'd11,  13'd186,  -13'd422,  13'd222,  13'd92,  -13'd419,  -13'd428,  -13'd297,  -13'd130,  -13'd324,  13'd525,  -13'd134,  13'd433,  13'd106,  13'd380,  13'd424,  
-13'd56,  -13'd252,  13'd350,  -13'd153,  -13'd326,  -13'd121,  -13'd60,  -13'd2,  -13'd508,  13'd333,  -13'd925,  -13'd497,  13'd159,  13'd77,  13'd475,  -13'd291,  
-13'd269,  13'd17,  13'd246,  -13'd213,  -13'd391,  -13'd417,  13'd378,  13'd72,  13'd131,  13'd193,  13'd103,  13'd164,  -13'd795,  13'd357,  -13'd230,  -13'd216,  
13'd604,  13'd949,  -13'd61,  -13'd98,  13'd441,  -13'd188,  -13'd364,  -13'd335,  -13'd1064,  13'd84,  13'd67,  -13'd105,  -13'd781,  13'd341,  -13'd439,  -13'd371,  
-13'd580,  13'd842,  13'd552,  13'd497,  13'd745,  13'd39,  -13'd241,  -13'd114,  13'd555,  13'd978,  -13'd219,  -13'd563,  13'd39,  -13'd168,  13'd732,  -13'd253,  
13'd19,  -13'd230,  -13'd434,  13'd227,  13'd592,  13'd298,  13'd206,  13'd557,  -13'd127,  13'd743,  13'd388,  13'd98,  -13'd548,  13'd85,  13'd356,  13'd737,  

-13'd1008,  -13'd17,  13'd78,  13'd148,  13'd180,  13'd306,  13'd42,  -13'd250,  13'd275,  13'd267,  13'd748,  -13'd709,  -13'd82,  -13'd228,  13'd1105,  -13'd115,  
-13'd555,  -13'd581,  -13'd761,  -13'd267,  13'd265,  -13'd382,  -13'd450,  13'd582,  13'd346,  13'd50,  13'd285,  -13'd257,  13'd181,  13'd181,  13'd12,  13'd205,  
13'd106,  -13'd1305,  13'd570,  13'd591,  13'd550,  -13'd549,  13'd55,  13'd350,  -13'd221,  -13'd119,  13'd195,  13'd493,  -13'd266,  -13'd613,  13'd510,  -13'd625,  
13'd111,  -13'd743,  13'd222,  13'd285,  -13'd466,  13'd408,  13'd330,  -13'd92,  13'd367,  -13'd127,  13'd281,  13'd206,  -13'd398,  -13'd26,  -13'd212,  -13'd367,  
-13'd842,  -13'd493,  13'd429,  -13'd260,  -13'd428,  13'd122,  -13'd161,  13'd565,  -13'd372,  13'd457,  -13'd406,  -13'd368,  -13'd90,  -13'd120,  -13'd182,  -13'd653,  
13'd145,  13'd361,  13'd142,  -13'd436,  -13'd351,  -13'd358,  -13'd875,  13'd284,  -13'd662,  13'd284,  13'd159,  13'd567,  -13'd459,  13'd423,  -13'd580,  -13'd763,  
-13'd381,  -13'd353,  -13'd933,  -13'd465,  13'd383,  13'd303,  13'd341,  -13'd915,  -13'd348,  -13'd348,  13'd308,  13'd164,  -13'd324,  -13'd342,  13'd144,  -13'd287,  
-13'd3,  13'd91,  13'd14,  13'd452,  -13'd28,  13'd522,  -13'd700,  13'd170,  -13'd684,  13'd37,  -13'd59,  13'd499,  -13'd177,  -13'd65,  -13'd383,  13'd797,  
-13'd567,  13'd261,  -13'd316,  13'd1005,  13'd530,  13'd595,  13'd713,  -13'd397,  -13'd397,  -13'd1,  13'd293,  -13'd238,  -13'd18,  13'd1135,  13'd272,  13'd351,  
-13'd823,  -13'd1225,  -13'd156,  -13'd706,  13'd255,  -13'd451,  13'd346,  13'd395,  -13'd474,  13'd204,  -13'd243,  -13'd732,  -13'd682,  13'd462,  -13'd437,  13'd108,  
13'd211,  13'd553,  13'd364,  13'd79,  -13'd203,  -13'd202,  -13'd7,  13'd531,  -13'd232,  -13'd711,  13'd731,  13'd192,  -13'd776,  13'd520,  -13'd610,  -13'd480,  
13'd183,  -13'd8,  -13'd826,  -13'd713,  13'd153,  -13'd560,  13'd718,  -13'd226,  -13'd339,  13'd439,  -13'd32,  13'd643,  13'd95,  13'd243,  13'd604,  13'd638,  
13'd307,  13'd384,  13'd412,  13'd701,  -13'd210,  13'd268,  13'd143,  13'd354,  -13'd83,  13'd362,  13'd259,  13'd617,  13'd572,  13'd152,  13'd87,  -13'd37,  
13'd105,  -13'd263,  13'd461,  13'd156,  13'd33,  13'd499,  13'd490,  -13'd387,  -13'd21,  -13'd1261,  13'd75,  13'd362,  -13'd512,  -13'd183,  13'd637,  -13'd41,  
-13'd738,  -13'd696,  13'd940,  13'd423,  13'd161,  13'd260,  13'd28,  -13'd401,  -13'd746,  -13'd70,  -13'd148,  13'd492,  -13'd284,  -13'd126,  -13'd472,  -13'd402,  
-13'd200,  13'd281,  13'd536,  -13'd819,  -13'd719,  13'd193,  13'd686,  -13'd248,  -13'd366,  -13'd61,  13'd337,  13'd132,  -13'd315,  13'd285,  -13'd179,  13'd429,  
-13'd24,  13'd214,  -13'd195,  -13'd474,  13'd6,  -13'd247,  13'd765,  -13'd248,  13'd291,  -13'd379,  13'd189,  13'd61,  13'd370,  -13'd250,  13'd223,  13'd62,  
13'd176,  13'd57,  13'd486,  13'd369,  -13'd488,  -13'd89,  13'd163,  13'd739,  13'd36,  -13'd360,  13'd175,  -13'd181,  13'd11,  13'd127,  -13'd206,  13'd55,  
13'd302,  13'd233,  13'd549,  -13'd50,  -13'd481,  -13'd138,  13'd657,  13'd635,  13'd595,  -13'd1181,  13'd920,  -13'd180,  13'd624,  -13'd904,  -13'd382,  -13'd131,  
13'd588,  13'd239,  -13'd249,  -13'd374,  -13'd297,  -13'd28,  -13'd204,  13'd608,  -13'd908,  -13'd1410,  -13'd36,  13'd64,  13'd427,  13'd592,  13'd902,  13'd444,  
-13'd141,  -13'd791,  -13'd641,  -13'd692,  -13'd434,  -13'd871,  13'd865,  13'd115,  -13'd528,  13'd462,  13'd138,  -13'd410,  -13'd279,  13'd67,  13'd103,  -13'd59,  
-13'd265,  13'd156,  13'd508,  -13'd119,  -13'd78,  13'd521,  13'd1240,  13'd526,  13'd267,  13'd566,  -13'd225,  13'd194,  13'd285,  13'd524,  -13'd355,  -13'd243,  
-13'd347,  13'd535,  13'd950,  -13'd994,  13'd675,  -13'd1276,  13'd246,  13'd382,  13'd611,  -13'd110,  -13'd412,  -13'd867,  -13'd498,  13'd263,  13'd682,  -13'd510,  
13'd90,  -13'd382,  -13'd392,  -13'd190,  -13'd443,  -13'd951,  -13'd23,  13'd207,  -13'd301,  -13'd841,  -13'd721,  -13'd1075,  -13'd1015,  -13'd79,  -13'd689,  -13'd186,  
-13'd347,  -13'd293,  13'd493,  -13'd508,  -13'd975,  -13'd396,  -13'd17,  13'd269,  -13'd395,  -13'd564,  -13'd540,  -13'd669,  -13'd628,  -13'd624,  -13'd411,  -13'd777,  

-13'd254,  -13'd466,  13'd190,  13'd101,  13'd67,  -13'd77,  -13'd822,  13'd837,  13'd66,  13'd534,  -13'd221,  -13'd363,  -13'd160,  -13'd118,  13'd903,  13'd784,  
-13'd260,  -13'd654,  13'd186,  13'd434,  13'd89,  13'd202,  -13'd803,  13'd280,  -13'd449,  13'd714,  13'd782,  13'd108,  13'd673,  -13'd480,  13'd439,  13'd160,  
13'd425,  -13'd10,  -13'd170,  13'd268,  13'd99,  13'd127,  13'd61,  -13'd330,  -13'd812,  13'd52,  13'd409,  13'd79,  13'd332,  -13'd1840,  -13'd697,  13'd554,  
13'd774,  -13'd22,  -13'd156,  13'd109,  -13'd157,  13'd713,  13'd416,  -13'd125,  13'd663,  -13'd366,  13'd337,  13'd435,  -13'd203,  -13'd710,  -13'd209,  -13'd84,  
13'd542,  -13'd708,  13'd748,  -13'd147,  -13'd1,  -13'd203,  13'd322,  -13'd294,  13'd191,  13'd278,  -13'd295,  -13'd28,  -13'd587,  -13'd163,  -13'd471,  13'd223,  
-13'd256,  13'd324,  -13'd143,  -13'd98,  13'd573,  13'd432,  -13'd524,  13'd371,  13'd591,  -13'd185,  13'd229,  13'd367,  13'd705,  13'd11,  13'd30,  -13'd540,  
-13'd531,  -13'd450,  -13'd884,  13'd715,  13'd204,  -13'd389,  -13'd825,  -13'd275,  -13'd615,  -13'd185,  13'd290,  13'd416,  13'd662,  -13'd266,  13'd230,  -13'd288,  
13'd525,  -13'd337,  -13'd694,  13'd634,  13'd519,  13'd200,  -13'd718,  13'd572,  -13'd319,  13'd154,  13'd107,  13'd68,  13'd217,  -13'd215,  13'd175,  13'd520,  
13'd372,  13'd168,  -13'd703,  13'd200,  13'd322,  13'd105,  13'd734,  13'd735,  13'd443,  13'd396,  13'd890,  -13'd367,  13'd314,  13'd45,  -13'd72,  13'd277,  
13'd91,  -13'd1118,  -13'd320,  13'd182,  -13'd525,  13'd211,  -13'd541,  13'd565,  13'd401,  13'd551,  13'd161,  -13'd190,  13'd539,  -13'd64,  -13'd181,  -13'd252,  
-13'd527,  13'd641,  -13'd224,  13'd489,  13'd553,  -13'd351,  13'd107,  13'd229,  13'd1250,  13'd269,  13'd633,  13'd200,  -13'd27,  13'd465,  -13'd2,  13'd43,  
-13'd437,  -13'd100,  -13'd234,  13'd294,  13'd24,  -13'd902,  -13'd874,  -13'd392,  -13'd710,  -13'd121,  13'd555,  -13'd48,  13'd660,  -13'd224,  -13'd43,  13'd402,  
-13'd7,  -13'd323,  13'd622,  13'd154,  -13'd793,  13'd706,  13'd462,  13'd110,  -13'd464,  13'd946,  13'd314,  13'd429,  13'd306,  -13'd726,  -13'd351,  13'd663,  
13'd219,  13'd343,  -13'd676,  13'd1,  13'd364,  13'd775,  -13'd174,  13'd605,  -13'd183,  -13'd324,  -13'd148,  13'd301,  13'd75,  13'd96,  13'd276,  13'd153,  
-13'd665,  -13'd281,  -13'd414,  -13'd16,  13'd702,  -13'd338,  -13'd320,  -13'd54,  13'd150,  -13'd98,  13'd543,  13'd227,  13'd730,  13'd26,  13'd397,  -13'd613,  
-13'd149,  13'd153,  -13'd576,  -13'd690,  13'd262,  -13'd101,  -13'd364,  13'd130,  13'd554,  -13'd19,  13'd320,  13'd192,  -13'd190,  -13'd542,  -13'd895,  -13'd401,  
-13'd1000,  -13'd690,  13'd350,  13'd290,  -13'd409,  -13'd471,  -13'd240,  -13'd739,  13'd73,  13'd339,  -13'd7,  13'd79,  -13'd495,  -13'd716,  13'd105,  13'd780,  
-13'd747,  13'd131,  -13'd33,  13'd123,  13'd160,  -13'd211,  13'd75,  -13'd405,  13'd887,  -13'd2,  13'd113,  13'd122,  13'd265,  -13'd914,  -13'd225,  -13'd291,  
-13'd136,  13'd360,  13'd343,  -13'd707,  -13'd569,  13'd444,  -13'd50,  -13'd240,  -13'd230,  13'd381,  13'd22,  13'd153,  -13'd2,  -13'd596,  -13'd647,  -13'd195,  
13'd447,  -13'd288,  -13'd335,  13'd192,  -13'd108,  -13'd203,  -13'd443,  13'd1003,  -13'd422,  13'd316,  -13'd130,  13'd84,  13'd445,  13'd329,  -13'd147,  13'd259,  
13'd368,  13'd565,  -13'd376,  -13'd213,  13'd741,  13'd429,  13'd625,  -13'd893,  13'd476,  13'd502,  -13'd113,  13'd63,  13'd164,  -13'd452,  -13'd601,  13'd149,  
-13'd200,  -13'd333,  13'd165,  -13'd715,  -13'd206,  13'd524,  13'd585,  -13'd125,  13'd424,  13'd835,  -13'd383,  -13'd442,  -13'd224,  13'd496,  -13'd237,  13'd403,  
13'd63,  13'd823,  13'd433,  -13'd83,  -13'd278,  13'd28,  13'd918,  -13'd187,  13'd244,  13'd565,  -13'd218,  -13'd424,  13'd218,  -13'd354,  13'd381,  13'd10,  
13'd47,  -13'd621,  13'd63,  -13'd346,  13'd205,  13'd79,  13'd45,  -13'd136,  13'd401,  -13'd347,  -13'd637,  -13'd1065,  -13'd1115,  13'd570,  13'd73,  13'd237,  
13'd245,  -13'd269,  13'd534,  -13'd596,  -13'd211,  -13'd326,  -13'd384,  -13'd442,  13'd317,  -13'd418,  -13'd150,  -13'd217,  13'd204,  -13'd624,  -13'd561,  13'd38,  

13'd795,  13'd85,  13'd70,  -13'd29,  -13'd230,  -13'd483,  13'd385,  13'd17,  13'd211,  -13'd232,  -13'd275,  -13'd294,  13'd11,  13'd74,  -13'd946,  -13'd408,  
13'd1120,  13'd155,  13'd542,  -13'd128,  -13'd19,  13'd306,  13'd647,  -13'd33,  13'd103,  -13'd53,  13'd431,  13'd265,  13'd40,  13'd201,  -13'd247,  13'd803,  
13'd957,  13'd55,  13'd74,  13'd617,  -13'd161,  -13'd592,  13'd185,  13'd278,  -13'd198,  -13'd125,  13'd410,  13'd45,  13'd758,  -13'd455,  13'd152,  13'd183,  
-13'd435,  13'd420,  13'd790,  13'd158,  -13'd68,  13'd497,  -13'd1225,  -13'd434,  -13'd817,  -13'd205,  -13'd288,  -13'd506,  13'd377,  -13'd280,  13'd89,  -13'd272,  
13'd226,  -13'd206,  13'd100,  -13'd24,  13'd836,  -13'd625,  -13'd219,  -13'd551,  -13'd1068,  -13'd383,  -13'd125,  -13'd558,  13'd661,  13'd192,  13'd10,  13'd1266,  
13'd646,  -13'd845,  13'd759,  -13'd127,  -13'd26,  13'd704,  -13'd156,  13'd499,  -13'd20,  -13'd85,  -13'd623,  -13'd426,  13'd34,  13'd274,  13'd102,  -13'd516,  
-13'd107,  -13'd507,  -13'd67,  -13'd273,  -13'd138,  -13'd51,  -13'd167,  -13'd235,  -13'd436,  13'd20,  13'd190,  13'd618,  -13'd500,  -13'd337,  -13'd14,  -13'd317,  
-13'd147,  13'd226,  -13'd416,  -13'd452,  13'd641,  13'd383,  13'd33,  13'd175,  13'd503,  13'd900,  13'd574,  -13'd66,  -13'd176,  -13'd309,  -13'd136,  13'd161,  
-13'd190,  -13'd40,  -13'd144,  -13'd189,  13'd242,  -13'd544,  -13'd928,  13'd188,  -13'd420,  13'd1034,  13'd535,  -13'd161,  13'd111,  -13'd662,  -13'd542,  13'd397,  
-13'd288,  -13'd99,  -13'd309,  -13'd282,  13'd931,  13'd475,  -13'd444,  13'd338,  -13'd186,  13'd290,  13'd186,  13'd91,  -13'd45,  13'd94,  -13'd376,  13'd384,  
13'd105,  13'd18,  13'd89,  -13'd265,  13'd428,  -13'd6,  -13'd453,  -13'd219,  -13'd558,  13'd288,  -13'd639,  13'd215,  -13'd628,  13'd182,  13'd706,  -13'd215,  
-13'd337,  13'd130,  -13'd274,  13'd115,  13'd508,  13'd483,  -13'd340,  -13'd456,  13'd110,  13'd142,  13'd32,  13'd30,  -13'd361,  -13'd558,  13'd74,  -13'd93,  
13'd150,  -13'd414,  13'd151,  13'd663,  13'd459,  13'd53,  -13'd48,  13'd639,  13'd957,  -13'd94,  -13'd103,  13'd220,  -13'd968,  -13'd226,  -13'd177,  13'd23,  
13'd712,  -13'd318,  -13'd316,  -13'd186,  -13'd274,  13'd196,  -13'd331,  -13'd92,  13'd451,  13'd1288,  13'd89,  -13'd303,  13'd468,  13'd218,  -13'd1056,  13'd133,  
13'd305,  13'd299,  -13'd604,  -13'd221,  13'd794,  13'd335,  -13'd169,  -13'd483,  13'd243,  13'd806,  13'd326,  13'd469,  -13'd399,  -13'd2,  -13'd426,  -13'd120,  
13'd496,  13'd235,  -13'd209,  13'd536,  -13'd63,  -13'd683,  13'd212,  -13'd126,  -13'd486,  13'd438,  -13'd731,  13'd299,  13'd37,  13'd374,  13'd202,  13'd255,  
13'd798,  13'd738,  13'd279,  13'd830,  -13'd22,  -13'd159,  13'd36,  -13'd304,  13'd700,  13'd715,  -13'd63,  13'd542,  -13'd238,  13'd340,  13'd233,  -13'd617,  
13'd518,  13'd638,  -13'd35,  13'd198,  13'd698,  13'd118,  -13'd591,  -13'd179,  -13'd346,  -13'd233,  13'd487,  13'd173,  -13'd275,  13'd426,  -13'd108,  13'd416,  
-13'd389,  13'd424,  -13'd513,  -13'd173,  13'd310,  -13'd751,  -13'd492,  13'd108,  -13'd475,  -13'd187,  -13'd110,  -13'd81,  13'd115,  -13'd172,  13'd1005,  -13'd356,  
13'd8,  -13'd225,  13'd365,  -13'd89,  -13'd834,  13'd681,  -13'd688,  13'd592,  13'd245,  13'd43,  -13'd25,  13'd525,  13'd559,  13'd413,  -13'd56,  13'd144,  
13'd616,  13'd35,  13'd150,  13'd367,  -13'd619,  13'd384,  13'd0,  13'd616,  13'd465,  13'd615,  -13'd14,  13'd347,  13'd14,  13'd1186,  -13'd22,  -13'd237,  
13'd165,  13'd113,  13'd71,  13'd586,  13'd452,  13'd45,  -13'd390,  13'd480,  13'd112,  -13'd206,  13'd405,  -13'd305,  13'd339,  13'd428,  13'd1008,  -13'd99,  
-13'd333,  -13'd217,  -13'd687,  13'd25,  13'd501,  13'd299,  -13'd340,  13'd125,  -13'd285,  -13'd686,  -13'd111,  -13'd96,  13'd460,  -13'd1327,  13'd261,  -13'd53,  
13'd305,  13'd117,  13'd177,  -13'd115,  13'd162,  13'd648,  13'd35,  13'd880,  13'd99,  -13'd164,  -13'd210,  13'd645,  13'd335,  13'd98,  -13'd38,  13'd281,  
13'd166,  13'd435,  13'd624,  -13'd1,  -13'd403,  13'd154,  13'd479,  13'd338,  13'd691,  13'd227,  -13'd565,  13'd1102,  -13'd429,  -13'd223,  13'd5,  13'd4,  

-13'd494,  13'd405,  -13'd322,  13'd231,  13'd893,  -13'd119,  -13'd713,  13'd396,  -13'd507,  13'd162,  -13'd100,  13'd115,  -13'd83,  13'd442,  -13'd115,  13'd1030,  
-13'd563,  13'd403,  13'd166,  13'd504,  13'd331,  13'd445,  -13'd347,  -13'd93,  13'd246,  13'd499,  -13'd697,  13'd385,  -13'd169,  -13'd782,  13'd927,  13'd1197,  
-13'd476,  -13'd70,  13'd558,  13'd258,  -13'd144,  -13'd458,  13'd93,  13'd286,  13'd31,  13'd36,  -13'd504,  13'd176,  13'd364,  13'd434,  -13'd611,  13'd607,  
-13'd253,  -13'd846,  13'd63,  -13'd9,  13'd89,  -13'd248,  13'd707,  -13'd403,  -13'd11,  -13'd324,  13'd282,  13'd593,  -13'd576,  13'd1363,  13'd68,  -13'd852,  
-13'd744,  13'd311,  13'd548,  -13'd564,  -13'd575,  -13'd245,  13'd168,  -13'd619,  13'd139,  -13'd165,  -13'd750,  -13'd562,  -13'd810,  13'd608,  -13'd750,  -13'd553,  
13'd496,  13'd618,  -13'd417,  -13'd332,  13'd344,  -13'd164,  -13'd253,  13'd339,  -13'd165,  -13'd570,  13'd175,  13'd24,  13'd196,  -13'd559,  13'd407,  13'd557,  
13'd73,  13'd240,  -13'd392,  -13'd455,  13'd144,  13'd335,  -13'd213,  -13'd306,  13'd83,  13'd1023,  13'd398,  13'd587,  -13'd165,  13'd15,  13'd537,  13'd188,  
13'd949,  13'd283,  13'd967,  13'd352,  -13'd537,  -13'd377,  13'd45,  -13'd24,  13'd94,  13'd279,  -13'd136,  13'd644,  13'd76,  -13'd448,  13'd86,  13'd11,  
13'd774,  -13'd396,  13'd319,  13'd678,  13'd31,  13'd758,  13'd891,  -13'd119,  -13'd526,  13'd396,  13'd167,  13'd274,  13'd79,  13'd1472,  -13'd272,  -13'd265,  
13'd457,  -13'd155,  13'd134,  13'd210,  13'd612,  13'd728,  13'd107,  -13'd831,  -13'd1,  -13'd563,  13'd200,  -13'd266,  13'd239,  13'd883,  -13'd907,  -13'd663,  
-13'd1094,  -13'd225,  -13'd517,  13'd16,  13'd12,  -13'd484,  13'd399,  13'd199,  13'd682,  13'd260,  -13'd136,  -13'd396,  -13'd245,  -13'd327,  -13'd886,  13'd285,  
13'd335,  13'd63,  -13'd15,  13'd25,  -13'd182,  -13'd139,  -13'd663,  13'd634,  -13'd482,  13'd3,  -13'd178,  -13'd352,  13'd375,  13'd749,  13'd315,  13'd11,  
13'd352,  -13'd422,  -13'd487,  -13'd96,  13'd57,  -13'd177,  -13'd101,  13'd575,  -13'd1374,  13'd212,  13'd449,  -13'd177,  13'd703,  -13'd173,  13'd384,  -13'd491,  
-13'd1,  -13'd301,  13'd448,  13'd769,  13'd200,  13'd338,  -13'd133,  13'd395,  -13'd233,  13'd235,  13'd637,  13'd231,  13'd395,  -13'd283,  -13'd470,  13'd94,  
-13'd299,  -13'd789,  -13'd55,  -13'd709,  13'd498,  13'd124,  -13'd62,  13'd251,  -13'd68,  13'd187,  13'd267,  13'd200,  13'd736,  13'd63,  -13'd546,  -13'd101,  
-13'd1189,  -13'd999,  13'd183,  13'd420,  13'd416,  -13'd1,  -13'd759,  13'd589,  13'd592,  -13'd57,  13'd25,  -13'd1036,  -13'd355,  -13'd103,  -13'd222,  -13'd490,  
-13'd592,  13'd91,  13'd331,  -13'd254,  13'd208,  13'd139,  -13'd371,  -13'd542,  -13'd147,  13'd318,  13'd195,  -13'd479,  -13'd297,  -13'd708,  -13'd45,  -13'd145,  
-13'd479,  13'd449,  13'd144,  -13'd324,  -13'd526,  -13'd310,  -13'd148,  13'd397,  13'd159,  13'd429,  13'd478,  13'd82,  -13'd672,  -13'd261,  13'd92,  13'd111,  
-13'd389,  -13'd118,  -13'd37,  -13'd668,  -13'd318,  13'd452,  -13'd363,  13'd167,  13'd214,  -13'd437,  13'd486,  -13'd303,  -13'd45,  13'd641,  -13'd366,  13'd92,  
13'd98,  13'd546,  13'd47,  -13'd548,  13'd204,  13'd48,  13'd100,  -13'd333,  -13'd135,  -13'd306,  13'd4,  -13'd410,  13'd475,  13'd46,  13'd115,  13'd223,  
-13'd609,  -13'd625,  -13'd162,  -13'd37,  13'd153,  -13'd168,  13'd1015,  -13'd446,  -13'd43,  -13'd22,  -13'd322,  13'd538,  13'd765,  -13'd405,  13'd425,  -13'd213,  
13'd944,  -13'd142,  13'd264,  -13'd275,  13'd619,  13'd114,  13'd503,  -13'd565,  13'd318,  -13'd107,  -13'd36,  13'd506,  -13'd358,  -13'd16,  13'd395,  13'd405,  
13'd397,  13'd803,  13'd290,  13'd24,  13'd116,  13'd199,  13'd95,  13'd117,  -13'd216,  -13'd421,  -13'd42,  13'd430,  13'd51,  13'd292,  -13'd474,  13'd156,  
-13'd245,  -13'd262,  13'd198,  -13'd391,  -13'd270,  -13'd664,  13'd588,  13'd54,  -13'd457,  13'd201,  13'd322,  13'd184,  -13'd73,  13'd484,  -13'd216,  13'd73,  
13'd384,  13'd428,  13'd447,  13'd423,  13'd369,  -13'd901,  13'd763,  -13'd294,  -13'd121,  13'd255,  13'd74,  13'd320,  -13'd328,  13'd375,  -13'd309,  -13'd374,  

-13'd105,  -13'd118,  -13'd257,  -13'd187,  -13'd608,  13'd189,  -13'd874,  -13'd37,  -13'd959,  -13'd331,  13'd980,  -13'd380,  -13'd4,  -13'd680,  13'd247,  13'd256,  
-13'd12,  13'd281,  -13'd869,  13'd363,  13'd728,  13'd598,  -13'd395,  13'd611,  13'd679,  -13'd107,  -13'd111,  13'd613,  13'd297,  -13'd711,  13'd295,  -13'd182,  
-13'd124,  13'd480,  13'd411,  -13'd143,  13'd333,  13'd410,  -13'd833,  13'd314,  13'd428,  -13'd610,  -13'd376,  13'd490,  13'd297,  -13'd907,  13'd267,  13'd303,  
13'd396,  -13'd156,  13'd792,  13'd74,  -13'd243,  13'd138,  13'd560,  13'd578,  13'd226,  13'd794,  13'd331,  -13'd121,  13'd972,  -13'd485,  13'd237,  13'd94,  
-13'd244,  -13'd1388,  -13'd229,  13'd79,  -13'd211,  13'd554,  13'd382,  -13'd229,  -13'd200,  13'd626,  13'd484,  -13'd508,  -13'd294,  -13'd449,  13'd42,  -13'd219,  
-13'd341,  -13'd603,  13'd11,  -13'd496,  13'd43,  -13'd168,  13'd127,  -13'd674,  -13'd349,  -13'd769,  13'd279,  -13'd432,  -13'd340,  13'd29,  -13'd414,  13'd179,  
13'd12,  13'd72,  -13'd853,  13'd98,  -13'd46,  13'd471,  13'd275,  -13'd454,  -13'd216,  13'd421,  -13'd120,  -13'd268,  13'd54,  -13'd84,  -13'd922,  13'd606,  
-13'd585,  13'd928,  -13'd346,  -13'd568,  -13'd121,  13'd78,  13'd130,  -13'd239,  13'd89,  13'd344,  13'd194,  -13'd409,  13'd130,  13'd970,  -13'd467,  -13'd221,  
13'd228,  13'd371,  13'd109,  -13'd122,  13'd23,  13'd835,  13'd731,  -13'd209,  13'd499,  -13'd335,  -13'd359,  13'd570,  -13'd35,  13'd1235,  13'd528,  13'd46,  
-13'd1211,  13'd919,  13'd677,  13'd188,  13'd222,  -13'd140,  -13'd401,  -13'd494,  -13'd81,  -13'd827,  13'd217,  -13'd835,  -13'd1085,  13'd376,  13'd1112,  -13'd467,  
-13'd627,  -13'd486,  -13'd505,  -13'd111,  -13'd491,  -13'd882,  13'd560,  -13'd519,  -13'd377,  13'd316,  13'd151,  13'd144,  -13'd537,  -13'd505,  13'd97,  -13'd389,  
-13'd52,  13'd50,  -13'd486,  13'd29,  -13'd41,  13'd123,  13'd313,  -13'd498,  13'd756,  -13'd55,  -13'd555,  13'd440,  13'd243,  -13'd1520,  -13'd153,  13'd186,  
-13'd162,  13'd110,  -13'd327,  -13'd722,  -13'd7,  -13'd645,  13'd460,  -13'd189,  13'd161,  13'd476,  -13'd51,  -13'd374,  -13'd116,  13'd346,  -13'd70,  -13'd30,  
13'd370,  13'd164,  13'd341,  13'd665,  -13'd321,  13'd172,  13'd171,  -13'd129,  13'd35,  -13'd968,  -13'd341,  13'd783,  -13'd283,  13'd114,  13'd273,  -13'd977,  
13'd940,  -13'd80,  -13'd184,  13'd672,  -13'd896,  13'd240,  -13'd176,  -13'd13,  -13'd98,  -13'd168,  -13'd45,  13'd528,  -13'd81,  13'd144,  13'd452,  -13'd801,  
13'd563,  -13'd545,  13'd481,  13'd457,  -13'd1380,  13'd41,  13'd737,  -13'd6,  13'd354,  13'd161,  13'd524,  13'd18,  -13'd271,  -13'd83,  -13'd51,  13'd299,  
13'd41,  -13'd857,  -13'd64,  -13'd180,  -13'd689,  -13'd152,  -13'd449,  -13'd9,  13'd243,  13'd311,  -13'd281,  13'd778,  13'd696,  -13'd287,  -13'd279,  13'd8,  
13'd555,  -13'd457,  13'd307,  -13'd108,  -13'd351,  13'd572,  -13'd308,  13'd434,  -13'd137,  -13'd247,  -13'd948,  13'd226,  13'd503,  13'd303,  13'd414,  -13'd105,  
13'd287,  13'd55,  13'd241,  13'd523,  -13'd81,  13'd343,  13'd374,  13'd596,  13'd844,  13'd696,  -13'd295,  13'd55,  -13'd46,  -13'd548,  -13'd355,  -13'd272,  
13'd553,  13'd368,  -13'd883,  13'd286,  -13'd30,  13'd362,  13'd77,  13'd378,  -13'd18,  13'd454,  13'd658,  13'd74,  13'd265,  13'd256,  13'd231,  13'd184,  
13'd165,  -13'd361,  13'd664,  -13'd471,  -13'd362,  13'd276,  -13'd10,  13'd76,  -13'd373,  -13'd72,  13'd159,  -13'd160,  -13'd91,  13'd412,  -13'd162,  13'd533,  
-13'd277,  13'd328,  -13'd701,  -13'd203,  -13'd81,  13'd531,  13'd424,  -13'd9,  13'd460,  -13'd680,  13'd515,  -13'd500,  13'd209,  13'd181,  13'd404,  13'd144,  
-13'd251,  13'd556,  13'd275,  -13'd188,  -13'd293,  -13'd362,  -13'd391,  13'd267,  -13'd494,  -13'd452,  13'd142,  -13'd438,  13'd358,  13'd611,  -13'd316,  -13'd402,  
-13'd816,  13'd300,  -13'd12,  13'd354,  -13'd80,  13'd230,  -13'd166,  13'd235,  -13'd419,  -13'd102,  -13'd22,  -13'd550,  13'd49,  13'd189,  13'd121,  13'd117,  
-13'd137,  -13'd345,  -13'd1018,  -13'd353,  -13'd215,  13'd243,  13'd300,  13'd149,  -13'd1161,  13'd1679,  13'd320,  13'd150,  -13'd320,  -13'd224,  -13'd352,  13'd566,  

-13'd369,  -13'd253,  13'd314,  -13'd468,  -13'd69,  -13'd364,  13'd1645,  -13'd464,  13'd604,  13'd200,  13'd298,  13'd74,  -13'd71,  13'd282,  13'd601,  13'd811,  
-13'd691,  13'd236,  13'd398,  -13'd709,  -13'd944,  13'd260,  13'd1456,  13'd60,  -13'd672,  13'd44,  13'd355,  13'd391,  13'd555,  13'd864,  -13'd314,  -13'd101,  
13'd327,  -13'd226,  13'd517,  -13'd917,  -13'd111,  -13'd351,  13'd910,  -13'd21,  -13'd724,  -13'd903,  13'd313,  13'd549,  -13'd868,  13'd955,  -13'd282,  -13'd1428,  
13'd1488,  13'd266,  -13'd790,  -13'd505,  -13'd171,  13'd42,  13'd726,  -13'd259,  -13'd519,  -13'd592,  -13'd25,  13'd172,  13'd89,  13'd514,  -13'd783,  -13'd620,  
13'd410,  13'd701,  -13'd233,  -13'd51,  -13'd877,  -13'd240,  13'd56,  -13'd354,  13'd201,  13'd29,  -13'd263,  -13'd349,  -13'd740,  -13'd24,  13'd102,  13'd146,  
13'd511,  -13'd335,  13'd508,  -13'd31,  13'd83,  -13'd688,  13'd1267,  -13'd583,  -13'd192,  13'd383,  13'd875,  -13'd369,  13'd80,  -13'd368,  13'd226,  13'd567,  
-13'd512,  13'd291,  13'd48,  -13'd122,  13'd523,  -13'd300,  13'd685,  -13'd736,  -13'd446,  -13'd357,  13'd620,  13'd77,  13'd184,  -13'd232,  -13'd1098,  -13'd181,  
13'd979,  13'd577,  13'd448,  -13'd528,  -13'd835,  13'd0,  -13'd535,  -13'd199,  -13'd162,  13'd245,  -13'd403,  13'd28,  13'd522,  13'd234,  13'd172,  13'd68,  
13'd808,  13'd923,  -13'd291,  13'd333,  -13'd177,  13'd692,  -13'd419,  -13'd424,  13'd551,  13'd428,  13'd143,  13'd276,  13'd174,  13'd268,  13'd69,  13'd47,  
-13'd9,  -13'd646,  13'd207,  13'd465,  13'd378,  -13'd837,  -13'd154,  -13'd67,  -13'd3,  -13'd15,  13'd73,  13'd652,  13'd522,  -13'd660,  13'd462,  13'd172,  
13'd109,  -13'd733,  -13'd14,  -13'd131,  -13'd215,  -13'd486,  13'd1405,  -13'd216,  -13'd254,  -13'd396,  13'd148,  13'd634,  -13'd1038,  -13'd1105,  13'd469,  -13'd660,  
13'd727,  -13'd710,  -13'd519,  -13'd313,  -13'd278,  13'd556,  -13'd564,  -13'd211,  13'd483,  -13'd692,  13'd198,  13'd101,  -13'd522,  -13'd80,  -13'd91,  13'd83,  
13'd760,  13'd282,  -13'd27,  -13'd217,  -13'd120,  -13'd464,  -13'd6,  -13'd101,  -13'd123,  -13'd111,  -13'd977,  -13'd294,  13'd356,  -13'd593,  -13'd189,  -13'd288,  
-13'd16,  13'd501,  -13'd401,  -13'd413,  -13'd88,  13'd672,  13'd162,  -13'd491,  13'd322,  13'd615,  -13'd164,  13'd256,  -13'd55,  13'd39,  -13'd101,  -13'd181,  
-13'd288,  -13'd91,  13'd353,  13'd714,  -13'd318,  13'd143,  -13'd46,  -13'd62,  -13'd362,  13'd241,  -13'd765,  13'd396,  13'd373,  -13'd29,  13'd444,  13'd0,  
13'd239,  13'd147,  13'd272,  13'd112,  13'd371,  13'd266,  13'd677,  13'd486,  -13'd59,  13'd138,  -13'd436,  13'd294,  -13'd95,  13'd119,  -13'd73,  13'd11,  
13'd12,  -13'd362,  13'd162,  13'd658,  13'd80,  -13'd340,  13'd120,  -13'd689,  13'd177,  13'd68,  13'd336,  -13'd303,  13'd206,  13'd420,  -13'd20,  13'd268,  
13'd339,  -13'd501,  13'd41,  13'd284,  -13'd882,  -13'd284,  -13'd520,  13'd695,  13'd464,  13'd690,  -13'd369,  -13'd345,  13'd783,  -13'd491,  13'd106,  -13'd3,  
13'd778,  -13'd576,  -13'd595,  13'd169,  -13'd741,  -13'd219,  -13'd498,  13'd366,  -13'd324,  -13'd193,  13'd716,  13'd95,  13'd943,  13'd451,  13'd223,  -13'd705,  
13'd119,  -13'd86,  13'd423,  13'd289,  -13'd27,  -13'd353,  13'd306,  13'd394,  13'd185,  13'd535,  -13'd394,  -13'd34,  13'd998,  -13'd199,  -13'd97,  13'd388,  
-13'd298,  13'd337,  13'd7,  13'd893,  13'd313,  13'd692,  -13'd485,  13'd190,  13'd631,  13'd251,  13'd351,  -13'd828,  -13'd144,  -13'd413,  -13'd136,  13'd247,  
13'd78,  -13'd410,  13'd14,  13'd195,  -13'd201,  -13'd686,  13'd551,  -13'd311,  13'd244,  13'd457,  13'd72,  -13'd650,  13'd473,  -13'd440,  -13'd374,  13'd99,  
-13'd295,  13'd64,  -13'd433,  13'd13,  -13'd481,  13'd253,  -13'd34,  -13'd268,  -13'd80,  13'd888,  -13'd181,  13'd61,  13'd491,  -13'd676,  13'd204,  13'd704,  
-13'd1168,  -13'd391,  -13'd409,  13'd181,  13'd98,  13'd537,  -13'd351,  -13'd735,  -13'd322,  13'd556,  -13'd391,  -13'd490,  -13'd342,  -13'd337,  -13'd813,  13'd441,  
-13'd288,  -13'd48,  -13'd185,  -13'd188,  13'd221,  -13'd524,  -13'd836,  13'd134,  -13'd209,  -13'd307,  13'd476,  -13'd615,  13'd78,  -13'd61,  -13'd141,  -13'd86,  

-13'd250,  -13'd918,  -13'd67,  13'd350,  13'd401,  -13'd82,  -13'd716,  13'd181,  -13'd156,  13'd116,  13'd399,  -13'd95,  -13'd169,  -13'd333,  -13'd236,  -13'd929,  
-13'd111,  -13'd362,  -13'd825,  13'd668,  -13'd192,  13'd430,  -13'd345,  13'd785,  13'd113,  13'd612,  -13'd2,  -13'd277,  -13'd330,  -13'd473,  13'd601,  -13'd535,  
-13'd233,  -13'd58,  13'd133,  13'd761,  -13'd504,  13'd221,  -13'd366,  -13'd135,  -13'd138,  13'd200,  -13'd399,  -13'd110,  13'd503,  13'd302,  13'd642,  13'd517,  
13'd11,  -13'd265,  13'd614,  13'd70,  -13'd134,  -13'd242,  -13'd5,  13'd631,  -13'd60,  13'd720,  13'd214,  -13'd671,  -13'd357,  -13'd1328,  13'd611,  13'd673,  
13'd232,  13'd231,  13'd760,  -13'd56,  13'd119,  13'd383,  -13'd696,  13'd586,  13'd264,  -13'd163,  -13'd735,  13'd384,  13'd402,  13'd303,  13'd643,  -13'd673,  
-13'd432,  -13'd368,  13'd5,  -13'd187,  13'd699,  13'd230,  -13'd575,  -13'd11,  13'd65,  13'd285,  -13'd439,  -13'd406,  13'd701,  13'd401,  -13'd824,  13'd321,  
13'd521,  13'd568,  13'd653,  -13'd39,  -13'd287,  13'd907,  -13'd190,  13'd61,  -13'd224,  13'd383,  13'd915,  -13'd569,  13'd127,  13'd203,  13'd306,  13'd96,  
-13'd844,  13'd968,  13'd174,  -13'd2,  13'd82,  13'd671,  13'd2,  -13'd291,  13'd144,  -13'd152,  -13'd344,  -13'd619,  -13'd485,  13'd453,  13'd582,  13'd341,  
-13'd1104,  13'd975,  13'd629,  13'd674,  13'd728,  13'd443,  -13'd1001,  13'd472,  -13'd16,  -13'd198,  13'd93,  -13'd579,  -13'd306,  -13'd383,  13'd328,  13'd166,  
13'd422,  13'd630,  13'd592,  13'd374,  -13'd367,  13'd876,  13'd548,  13'd230,  -13'd61,  -13'd207,  -13'd17,  -13'd132,  -13'd278,  13'd57,  13'd642,  13'd399,  
-13'd502,  -13'd317,  13'd180,  -13'd756,  -13'd252,  -13'd404,  -13'd753,  -13'd313,  -13'd131,  -13'd54,  -13'd407,  13'd209,  -13'd22,  -13'd255,  -13'd338,  -13'd152,  
13'd363,  -13'd384,  13'd159,  -13'd311,  13'd234,  13'd383,  13'd142,  -13'd68,  -13'd80,  -13'd240,  13'd497,  -13'd50,  -13'd500,  13'd631,  13'd458,  13'd499,  
13'd56,  13'd15,  -13'd183,  -13'd100,  13'd470,  13'd273,  13'd369,  13'd544,  -13'd235,  -13'd468,  -13'd303,  -13'd246,  -13'd146,  13'd116,  -13'd151,  -13'd229,  
-13'd76,  13'd650,  13'd175,  13'd183,  -13'd9,  -13'd215,  13'd97,  -13'd308,  13'd483,  -13'd3,  13'd254,  -13'd214,  -13'd227,  13'd471,  13'd875,  -13'd485,  
13'd1344,  13'd663,  13'd372,  -13'd275,  13'd232,  -13'd723,  -13'd296,  -13'd364,  -13'd128,  -13'd320,  -13'd842,  -13'd50,  13'd343,  -13'd112,  13'd246,  -13'd80,  
13'd775,  -13'd16,  13'd232,  13'd158,  13'd561,  -13'd365,  13'd153,  -13'd715,  13'd590,  13'd209,  -13'd332,  13'd445,  -13'd841,  13'd200,  -13'd73,  13'd27,  
13'd883,  -13'd387,  13'd28,  -13'd63,  -13'd673,  13'd290,  13'd1033,  -13'd297,  13'd591,  -13'd20,  13'd326,  13'd668,  13'd269,  13'd274,  -13'd355,  -13'd110,  
-13'd44,  -13'd638,  -13'd352,  -13'd25,  13'd677,  13'd437,  -13'd34,  -13'd162,  13'd117,  13'd521,  13'd554,  13'd12,  13'd338,  13'd858,  -13'd73,  -13'd6,  
-13'd433,  13'd62,  -13'd650,  13'd397,  13'd70,  -13'd826,  -13'd759,  -13'd327,  -13'd91,  13'd60,  -13'd669,  13'd270,  -13'd227,  -13'd497,  -13'd326,  -13'd794,  
13'd34,  -13'd73,  13'd714,  -13'd374,  13'd99,  -13'd417,  -13'd569,  -13'd361,  -13'd556,  -13'd349,  13'd386,  -13'd65,  -13'd2,  -13'd919,  -13'd192,  13'd150,  
-13'd45,  13'd75,  13'd212,  -13'd135,  13'd83,  13'd625,  -13'd658,  13'd625,  -13'd80,  -13'd31,  13'd125,  13'd119,  13'd225,  13'd555,  13'd68,  -13'd173,  
-13'd347,  13'd466,  13'd377,  13'd114,  -13'd170,  13'd201,  -13'd110,  -13'd81,  13'd269,  -13'd527,  13'd198,  13'd44,  -13'd109,  13'd789,  13'd665,  13'd258,  
13'd255,  -13'd599,  13'd530,  -13'd237,  13'd454,  13'd43,  -13'd550,  -13'd11,  -13'd332,  -13'd142,  13'd64,  -13'd32,  13'd130,  -13'd580,  13'd709,  13'd223,  
-13'd298,  -13'd462,  -13'd288,  -13'd58,  13'd125,  13'd222,  13'd105,  13'd235,  -13'd252,  -13'd785,  13'd768,  13'd434,  13'd553,  13'd250,  -13'd474,  -13'd55,  
13'd662,  -13'd178,  13'd384,  -13'd689,  -13'd637,  -13'd249,  13'd190,  13'd105,  13'd210,  -13'd841,  -13'd130,  13'd282,  -13'd469,  -13'd68,  -13'd821,  -13'd491,  

13'd82,  -13'd102,  13'd933,  -13'd186,  13'd78,  -13'd334,  13'd706,  -13'd461,  13'd489,  13'd236,  -13'd170,  -13'd308,  -13'd362,  13'd556,  -13'd279,  -13'd877,  
-13'd63,  -13'd447,  13'd19,  13'd275,  13'd120,  13'd345,  13'd1374,  13'd48,  13'd42,  -13'd567,  13'd106,  13'd186,  13'd186,  13'd74,  -13'd389,  -13'd568,  
13'd271,  13'd750,  -13'd407,  -13'd61,  13'd169,  -13'd214,  -13'd147,  -13'd80,  13'd632,  -13'd496,  13'd404,  -13'd232,  13'd641,  -13'd125,  -13'd883,  -13'd447,  
13'd242,  13'd840,  -13'd425,  13'd494,  -13'd414,  13'd750,  -13'd247,  -13'd324,  -13'd142,  -13'd496,  13'd40,  13'd419,  13'd694,  -13'd231,  13'd252,  13'd587,  
13'd575,  13'd831,  -13'd61,  13'd371,  -13'd131,  -13'd373,  -13'd303,  13'd375,  -13'd734,  -13'd138,  -13'd168,  -13'd387,  13'd1409,  13'd157,  13'd213,  13'd575,  
13'd516,  -13'd204,  13'd700,  13'd508,  -13'd315,  13'd50,  -13'd146,  13'd96,  13'd905,  13'd942,  -13'd694,  13'd65,  13'd1211,  13'd442,  13'd830,  -13'd173,  
-13'd380,  13'd363,  13'd323,  -13'd172,  13'd122,  -13'd401,  -13'd617,  -13'd242,  13'd10,  13'd152,  -13'd17,  -13'd75,  -13'd505,  -13'd7,  13'd661,  13'd41,  
13'd94,  -13'd69,  -13'd254,  -13'd549,  -13'd421,  -13'd537,  -13'd308,  -13'd485,  13'd476,  13'd497,  13'd1053,  -13'd387,  13'd5,  -13'd324,  -13'd79,  13'd203,  
-13'd697,  13'd57,  -13'd307,  -13'd267,  -13'd572,  13'd0,  -13'd206,  -13'd1184,  -13'd278,  13'd264,  -13'd199,  13'd42,  13'd537,  -13'd647,  -13'd474,  13'd283,  
13'd424,  -13'd556,  -13'd639,  -13'd274,  13'd330,  13'd420,  -13'd669,  13'd272,  -13'd350,  13'd944,  13'd179,  13'd331,  13'd326,  -13'd245,  13'd249,  13'd66,  
-13'd296,  13'd732,  13'd552,  13'd769,  13'd286,  13'd246,  -13'd1371,  -13'd429,  13'd4,  13'd236,  -13'd484,  -13'd132,  13'd74,  13'd966,  13'd616,  13'd94,  
-13'd204,  13'd395,  13'd3,  13'd317,  -13'd314,  -13'd73,  13'd137,  -13'd82,  -13'd407,  -13'd259,  13'd261,  13'd370,  -13'd234,  13'd600,  13'd101,  -13'd13,  
-13'd919,  -13'd654,  -13'd647,  -13'd13,  13'd424,  13'd467,  13'd279,  -13'd117,  13'd474,  -13'd1200,  -13'd158,  13'd523,  -13'd84,  -13'd717,  -13'd96,  -13'd543,  
-13'd460,  13'd503,  -13'd767,  13'd309,  13'd805,  -13'd791,  -13'd197,  13'd29,  13'd338,  13'd440,  13'd82,  13'd126,  13'd76,  13'd240,  -13'd305,  -13'd32,  
-13'd580,  -13'd588,  -13'd385,  13'd304,  13'd424,  13'd634,  -13'd1091,  -13'd40,  13'd98,  13'd1154,  13'd206,  13'd464,  13'd448,  13'd101,  -13'd10,  -13'd381,  
-13'd120,  -13'd126,  13'd626,  -13'd148,  13'd330,  13'd62,  13'd338,  13'd298,  -13'd227,  -13'd280,  -13'd417,  13'd206,  -13'd224,  13'd295,  -13'd206,  -13'd308,  
13'd583,  13'd54,  13'd569,  -13'd72,  -13'd174,  -13'd358,  -13'd459,  13'd620,  13'd239,  13'd523,  -13'd195,  13'd805,  -13'd162,  13'd719,  13'd583,  13'd125,  
-13'd299,  13'd155,  -13'd500,  -13'd162,  13'd627,  13'd579,  13'd6,  13'd306,  -13'd415,  -13'd308,  13'd56,  13'd516,  -13'd546,  -13'd1332,  13'd396,  13'd532,  
-13'd550,  -13'd186,  -13'd507,  -13'd717,  13'd718,  -13'd36,  -13'd433,  -13'd865,  13'd167,  -13'd163,  13'd446,  -13'd585,  13'd158,  13'd319,  13'd662,  13'd578,  
-13'd356,  -13'd459,  13'd1155,  -13'd194,  -13'd250,  -13'd113,  -13'd94,  -13'd562,  13'd317,  -13'd475,  -13'd5,  13'd180,  -13'd20,  13'd31,  -13'd826,  -13'd384,  
13'd504,  -13'd607,  -13'd1,  -13'd541,  13'd83,  13'd269,  -13'd51,  13'd434,  13'd867,  -13'd449,  -13'd464,  13'd17,  13'd38,  13'd784,  -13'd6,  13'd17,  
13'd660,  13'd255,  13'd124,  13'd364,  13'd349,  -13'd639,  -13'd659,  -13'd175,  -13'd105,  -13'd152,  -13'd178,  -13'd3,  13'd469,  -13'd6,  13'd700,  13'd255,  
-13'd39,  -13'd79,  -13'd547,  -13'd147,  -13'd226,  13'd311,  13'd252,  13'd187,  -13'd310,  -13'd1140,  -13'd22,  13'd13,  13'd299,  -13'd875,  13'd379,  13'd37,  
-13'd407,  -13'd494,  -13'd650,  -13'd720,  -13'd358,  13'd124,  -13'd260,  13'd526,  13'd523,  -13'd948,  13'd437,  13'd358,  13'd419,  13'd600,  -13'd258,  -13'd163,  
-13'd60,  13'd258,  -13'd1069,  -13'd122,  -13'd521,  13'd111,  13'd226,  13'd494,  -13'd189,  -13'd1853,  13'd57,  -13'd31,  -13'd272,  -13'd421,  -13'd120,  -13'd331,  

-13'd276,  13'd164,  13'd547,  -13'd156,  -13'd150,  13'd224,  13'd780,  -13'd151,  13'd319,  13'd500,  -13'd484,  13'd318,  13'd465,  13'd1176,  -13'd261,  13'd137,  
13'd383,  13'd223,  13'd521,  -13'd231,  -13'd305,  13'd516,  13'd671,  13'd353,  13'd208,  13'd113,  13'd308,  13'd442,  13'd693,  13'd349,  -13'd414,  13'd676,  
13'd4,  13'd207,  -13'd80,  13'd39,  -13'd184,  13'd76,  13'd330,  13'd411,  13'd412,  -13'd3,  -13'd185,  13'd289,  13'd187,  -13'd224,  13'd327,  13'd187,  
-13'd336,  -13'd155,  13'd41,  -13'd29,  13'd404,  -13'd280,  -13'd367,  -13'd65,  -13'd686,  -13'd491,  -13'd112,  -13'd652,  -13'd254,  -13'd648,  -13'd333,  -13'd386,  
-13'd558,  13'd1126,  13'd337,  13'd1,  -13'd155,  13'd426,  13'd69,  13'd44,  -13'd631,  -13'd618,  13'd95,  13'd628,  -13'd283,  13'd843,  13'd179,  13'd1023,  
-13'd367,  13'd345,  13'd225,  -13'd476,  13'd427,  13'd74,  -13'd256,  -13'd41,  13'd250,  13'd429,  -13'd402,  13'd30,  13'd869,  13'd477,  -13'd679,  -13'd136,  
13'd426,  -13'd248,  -13'd65,  -13'd104,  13'd664,  13'd65,  -13'd524,  -13'd220,  -13'd712,  13'd237,  -13'd218,  13'd128,  -13'd62,  13'd475,  -13'd93,  -13'd218,  
-13'd656,  13'd44,  13'd22,  -13'd178,  13'd121,  -13'd380,  -13'd279,  13'd177,  13'd155,  -13'd341,  13'd479,  13'd257,  -13'd374,  13'd548,  -13'd171,  13'd188,  
-13'd692,  -13'd313,  13'd240,  -13'd342,  -13'd12,  -13'd226,  -13'd66,  13'd745,  13'd363,  13'd244,  13'd139,  -13'd675,  -13'd198,  -13'd601,  13'd396,  -13'd213,  
-13'd508,  13'd292,  13'd117,  -13'd187,  13'd156,  13'd19,  -13'd332,  13'd13,  13'd272,  13'd1055,  13'd197,  13'd400,  13'd208,  -13'd316,  13'd340,  13'd699,  
13'd40,  13'd236,  -13'd677,  -13'd320,  13'd345,  13'd467,  13'd481,  13'd322,  -13'd559,  13'd527,  -13'd375,  13'd476,  -13'd935,  -13'd491,  13'd340,  13'd173,  
-13'd116,  13'd89,  13'd721,  -13'd90,  13'd333,  13'd173,  -13'd660,  -13'd662,  13'd62,  13'd376,  13'd115,  13'd668,  -13'd179,  -13'd325,  -13'd767,  13'd208,  
-13'd743,  13'd899,  13'd41,  13'd274,  13'd654,  13'd100,  13'd75,  13'd559,  13'd42,  13'd755,  13'd529,  13'd44,  -13'd261,  -13'd506,  -13'd396,  13'd180,  
-13'd722,  13'd291,  -13'd190,  -13'd52,  13'd21,  13'd418,  -13'd618,  -13'd1,  13'd169,  13'd497,  -13'd47,  -13'd262,  -13'd166,  -13'd361,  -13'd213,  13'd48,  
13'd207,  -13'd476,  -13'd43,  13'd462,  13'd207,  13'd45,  13'd45,  -13'd10,  13'd640,  -13'd257,  13'd115,  13'd1,  -13'd370,  13'd237,  -13'd624,  13'd838,  
13'd565,  13'd456,  13'd60,  13'd130,  -13'd334,  13'd447,  13'd632,  13'd641,  13'd232,  -13'd388,  13'd443,  13'd564,  13'd561,  13'd832,  13'd354,  13'd672,  
13'd326,  13'd476,  13'd295,  13'd54,  13'd168,  13'd472,  13'd266,  -13'd808,  13'd346,  13'd762,  -13'd120,  13'd226,  -13'd151,  13'd60,  13'd417,  13'd209,  
-13'd180,  13'd429,  -13'd740,  13'd176,  13'd265,  13'd314,  13'd96,  13'd1,  -13'd362,  -13'd152,  -13'd233,  -13'd96,  -13'd687,  -13'd742,  13'd713,  -13'd355,  
-13'd776,  13'd534,  13'd178,  -13'd557,  13'd745,  13'd72,  -13'd37,  13'd125,  13'd216,  -13'd144,  -13'd363,  13'd705,  -13'd529,  13'd249,  -13'd76,  -13'd499,  
13'd379,  13'd248,  13'd998,  13'd284,  -13'd133,  13'd820,  -13'd22,  13'd122,  13'd268,  13'd164,  13'd369,  13'd103,  13'd126,  13'd534,  -13'd40,  -13'd202,  
13'd540,  13'd57,  13'd66,  -13'd55,  -13'd777,  13'd703,  -13'd602,  13'd876,  13'd222,  13'd51,  -13'd336,  -13'd214,  13'd77,  13'd1309,  -13'd314,  -13'd106,  
-13'd50,  13'd54,  13'd194,  13'd788,  13'd263,  13'd112,  -13'd536,  13'd581,  -13'd378,  13'd133,  -13'd152,  -13'd131,  13'd483,  13'd37,  13'd500,  13'd15,  
13'd326,  -13'd352,  -13'd514,  13'd362,  13'd235,  13'd589,  13'd136,  13'd124,  -13'd316,  -13'd680,  13'd695,  13'd247,  13'd1001,  -13'd1156,  13'd117,  -13'd1,  
13'd542,  13'd81,  -13'd114,  -13'd369,  -13'd92,  -13'd290,  13'd386,  13'd321,  13'd641,  -13'd80,  13'd143,  13'd678,  -13'd142,  -13'd135,  -13'd87,  -13'd629,  
13'd549,  -13'd342,  13'd228,  13'd96,  -13'd618,  13'd214,  -13'd436,  -13'd570,  13'd393,  -13'd90,  13'd137,  13'd615,  13'd731,  13'd779,  -13'd884,  13'd439,  

13'd97,  -13'd82,  -13'd594,  13'd529,  13'd301,  -13'd214,  -13'd146,  13'd37,  -13'd456,  13'd674,  13'd330,  -13'd161,  -13'd48,  -13'd417,  13'd71,  13'd441,  
-13'd119,  -13'd846,  -13'd155,  13'd360,  13'd235,  13'd337,  -13'd537,  13'd616,  13'd345,  -13'd59,  -13'd765,  -13'd557,  13'd745,  -13'd456,  13'd187,  13'd31,  
-13'd808,  -13'd139,  13'd469,  -13'd289,  13'd551,  -13'd275,  -13'd22,  13'd360,  -13'd383,  13'd372,  13'd103,  13'd535,  -13'd287,  -13'd441,  13'd43,  -13'd649,  
-13'd837,  -13'd1404,  13'd482,  -13'd539,  -13'd172,  -13'd409,  13'd112,  -13'd321,  -13'd246,  -13'd267,  13'd536,  13'd42,  -13'd785,  13'd705,  13'd747,  -13'd607,  
13'd81,  13'd207,  13'd144,  13'd277,  -13'd1004,  13'd222,  -13'd80,  13'd292,  13'd100,  -13'd267,  -13'd247,  13'd121,  -13'd818,  13'd74,  13'd717,  -13'd416,  
-13'd216,  13'd367,  -13'd88,  -13'd135,  -13'd55,  -13'd520,  13'd8,  -13'd378,  13'd252,  -13'd1020,  13'd426,  13'd245,  13'd586,  -13'd707,  13'd360,  13'd498,  
-13'd227,  13'd1092,  13'd266,  13'd318,  13'd656,  -13'd107,  13'd71,  -13'd424,  -13'd629,  -13'd395,  -13'd342,  13'd203,  13'd61,  -13'd819,  13'd348,  13'd890,  
-13'd58,  -13'd317,  -13'd153,  13'd547,  13'd339,  -13'd539,  -13'd254,  13'd208,  13'd288,  13'd223,  -13'd648,  13'd630,  -13'd268,  13'd165,  13'd16,  13'd413,  
13'd220,  -13'd130,  13'd165,  13'd356,  -13'd70,  -13'd24,  -13'd86,  -13'd106,  13'd82,  -13'd164,  13'd643,  13'd389,  13'd25,  -13'd683,  13'd571,  -13'd926,  
13'd1089,  13'd423,  13'd484,  -13'd1,  13'd267,  13'd124,  13'd51,  -13'd493,  13'd184,  -13'd45,  -13'd272,  -13'd472,  13'd740,  13'd422,  13'd285,  -13'd96,  
13'd89,  13'd421,  -13'd0,  -13'd448,  -13'd1192,  13'd385,  13'd334,  13'd28,  13'd630,  13'd100,  13'd735,  -13'd529,  13'd325,  13'd167,  -13'd581,  -13'd74,  
13'd125,  13'd904,  -13'd61,  -13'd154,  13'd32,  13'd461,  -13'd117,  13'd552,  13'd254,  13'd489,  -13'd822,  13'd901,  13'd177,  13'd229,  -13'd84,  -13'd144,  
-13'd299,  13'd665,  13'd239,  -13'd237,  13'd213,  13'd236,  13'd13,  13'd832,  -13'd247,  13'd373,  -13'd521,  -13'd397,  13'd716,  -13'd154,  13'd286,  -13'd741,  
-13'd1416,  -13'd450,  -13'd222,  13'd80,  -13'd196,  13'd183,  -13'd906,  -13'd32,  13'd60,  -13'd218,  -13'd612,  13'd94,  13'd590,  -13'd1247,  13'd391,  13'd609,  
-13'd520,  -13'd779,  -13'd609,  -13'd187,  13'd221,  -13'd736,  13'd5,  13'd384,  13'd560,  -13'd150,  -13'd253,  -13'd240,  13'd184,  13'd599,  -13'd221,  -13'd26,  
13'd40,  -13'd451,  13'd836,  13'd726,  -13'd573,  13'd827,  13'd8,  13'd385,  13'd234,  13'd92,  13'd365,  -13'd485,  -13'd284,  13'd73,  13'd192,  -13'd790,  
13'd925,  13'd267,  -13'd414,  -13'd145,  -13'd296,  13'd35,  -13'd100,  13'd115,  -13'd290,  -13'd138,  -13'd137,  13'd312,  -13'd672,  -13'd429,  13'd333,  -13'd290,  
13'd159,  13'd865,  -13'd308,  -13'd196,  -13'd39,  13'd75,  -13'd261,  13'd300,  -13'd393,  -13'd375,  13'd458,  -13'd19,  -13'd428,  -13'd384,  13'd731,  -13'd796,  
-13'd208,  13'd266,  -13'd46,  13'd595,  13'd842,  13'd2,  -13'd415,  -13'd181,  13'd147,  -13'd359,  -13'd157,  13'd802,  -13'd126,  13'd44,  13'd50,  -13'd156,  
-13'd285,  -13'd356,  13'd236,  13'd728,  -13'd518,  -13'd16,  -13'd4,  13'd1,  13'd252,  -13'd444,  -13'd26,  13'd136,  -13'd622,  13'd750,  13'd74,  13'd136,  
-13'd13,  -13'd97,  -13'd481,  -13'd436,  -13'd200,  13'd368,  13'd552,  13'd112,  13'd319,  13'd620,  13'd248,  -13'd19,  13'd172,  13'd157,  -13'd111,  -13'd431,  
13'd482,  13'd335,  -13'd553,  -13'd520,  13'd179,  -13'd133,  -13'd1055,  -13'd106,  13'd241,  13'd333,  13'd289,  13'd60,  -13'd501,  -13'd865,  13'd152,  -13'd299,  
13'd200,  -13'd210,  -13'd562,  -13'd3,  13'd31,  13'd419,  -13'd230,  -13'd98,  -13'd16,  -13'd34,  13'd107,  13'd824,  13'd251,  -13'd722,  13'd449,  13'd19,  
13'd857,  -13'd24,  13'd879,  -13'd125,  -13'd418,  13'd80,  -13'd132,  13'd553,  13'd1171,  13'd197,  13'd9,  13'd9,  -13'd401,  -13'd203,  -13'd245,  13'd89,  
13'd246,  13'd1316,  13'd661,  13'd23,  -13'd502,  -13'd574,  13'd113,  -13'd232,  13'd746,  -13'd1266,  -13'd122,  13'd157,  -13'd86,  13'd528,  13'd105,  -13'd300,  

-13'd402,  -13'd194,  13'd84,  13'd44,  13'd215,  13'd203,  13'd415,  13'd169,  -13'd491,  13'd716,  -13'd127,  13'd492,  13'd94,  13'd23,  13'd379,  -13'd453,  
13'd521,  -13'd18,  -13'd617,  13'd721,  13'd1191,  13'd1141,  -13'd126,  13'd693,  13'd491,  13'd634,  -13'd25,  13'd340,  13'd237,  -13'd493,  -13'd184,  13'd46,  
13'd643,  -13'd181,  -13'd51,  13'd110,  -13'd414,  -13'd167,  13'd655,  13'd574,  -13'd40,  -13'd177,  -13'd568,  13'd324,  13'd454,  -13'd1117,  13'd399,  13'd391,  
13'd431,  13'd184,  -13'd88,  -13'd104,  13'd407,  13'd414,  13'd775,  -13'd165,  -13'd717,  -13'd541,  13'd599,  13'd493,  13'd1062,  13'd331,  13'd373,  13'd569,  
-13'd297,  13'd306,  13'd71,  -13'd86,  13'd342,  -13'd252,  13'd578,  -13'd155,  13'd148,  13'd543,  -13'd271,  13'd123,  -13'd522,  13'd234,  13'd552,  -13'd497,  
-13'd58,  13'd616,  13'd238,  13'd745,  -13'd204,  -13'd566,  -13'd360,  -13'd305,  -13'd430,  -13'd441,  13'd1125,  13'd86,  13'd86,  13'd757,  13'd345,  13'd124,  
13'd350,  13'd832,  -13'd182,  13'd305,  13'd1122,  -13'd378,  13'd134,  -13'd725,  13'd298,  -13'd255,  13'd234,  13'd373,  -13'd256,  -13'd1324,  -13'd606,  13'd352,  
13'd145,  13'd165,  -13'd200,  -13'd641,  13'd122,  -13'd614,  13'd463,  -13'd399,  13'd1211,  13'd413,  13'd443,  13'd651,  -13'd376,  -13'd267,  -13'd377,  13'd1156,  
13'd666,  13'd421,  13'd98,  13'd156,  -13'd292,  -13'd393,  13'd97,  -13'd430,  13'd478,  -13'd134,  13'd917,  -13'd406,  13'd471,  -13'd391,  13'd93,  -13'd22,  
-13'd339,  13'd712,  -13'd794,  13'd14,  -13'd708,  13'd441,  13'd28,  -13'd319,  13'd719,  -13'd779,  13'd426,  -13'd1031,  13'd48,  13'd902,  13'd148,  13'd257,  
13'd157,  13'd334,  13'd678,  13'd267,  -13'd1454,  13'd125,  13'd752,  13'd113,  13'd57,  -13'd343,  13'd474,  -13'd618,  -13'd32,  -13'd164,  -13'd206,  13'd575,  
13'd217,  13'd534,  -13'd666,  -13'd1074,  -13'd58,  13'd125,  -13'd153,  -13'd628,  -13'd255,  -13'd420,  -13'd371,  -13'd128,  -13'd976,  13'd547,  -13'd556,  13'd199,  
13'd262,  13'd654,  -13'd101,  -13'd586,  -13'd265,  -13'd270,  -13'd152,  13'd218,  -13'd380,  13'd598,  -13'd301,  -13'd764,  13'd252,  13'd1107,  13'd499,  -13'd603,  
-13'd6,  13'd196,  -13'd281,  -13'd167,  13'd829,  -13'd179,  -13'd250,  -13'd190,  -13'd379,  13'd240,  -13'd3,  -13'd76,  -13'd380,  13'd246,  13'd328,  -13'd373,  
-13'd842,  13'd204,  13'd6,  -13'd248,  13'd666,  13'd205,  -13'd215,  13'd307,  -13'd254,  13'd68,  -13'd613,  -13'd548,  -13'd544,  13'd822,  13'd787,  13'd530,  
13'd89,  -13'd1022,  13'd29,  -13'd900,  -13'd330,  -13'd13,  13'd219,  -13'd132,  13'd437,  13'd416,  -13'd37,  -13'd600,  -13'd42,  13'd258,  -13'd1028,  -13'd833,  
13'd223,  13'd625,  13'd597,  -13'd90,  -13'd864,  -13'd291,  13'd551,  -13'd211,  -13'd665,  13'd65,  -13'd293,  -13'd437,  -13'd210,  13'd289,  13'd217,  -13'd579,  
-13'd426,  -13'd443,  13'd259,  -13'd920,  13'd242,  13'd302,  13'd560,  13'd131,  13'd143,  -13'd206,  13'd292,  13'd179,  -13'd646,  13'd243,  -13'd411,  13'd539,  
-13'd1229,  -13'd357,  -13'd1179,  13'd496,  13'd756,  13'd535,  13'd41,  -13'd483,  13'd131,  -13'd914,  -13'd631,  -13'd115,  -13'd462,  -13'd249,  13'd476,  -13'd202,  
-13'd271,  13'd268,  13'd477,  -13'd110,  13'd207,  13'd500,  13'd404,  -13'd743,  13'd459,  -13'd366,  -13'd435,  13'd368,  -13'd665,  -13'd243,  13'd535,  -13'd237,  
-13'd716,  -13'd108,  13'd214,  13'd758,  13'd382,  13'd158,  13'd819,  13'd475,  13'd686,  13'd278,  -13'd626,  -13'd221,  13'd417,  13'd250,  13'd717,  -13'd384,  
13'd329,  13'd99,  13'd180,  13'd99,  -13'd204,  -13'd312,  -13'd716,  13'd85,  -13'd201,  13'd543,  -13'd488,  13'd406,  -13'd761,  -13'd890,  13'd33,  -13'd290,  
-13'd52,  -13'd206,  -13'd1,  -13'd542,  -13'd185,  13'd180,  -13'd427,  -13'd52,  -13'd254,  13'd891,  -13'd425,  13'd337,  -13'd475,  -13'd412,  -13'd266,  13'd266,  
13'd371,  13'd544,  13'd546,  -13'd423,  -13'd317,  13'd255,  -13'd191,  -13'd212,  13'd181,  13'd345,  -13'd719,  13'd79,  -13'd42,  13'd308,  -13'd156,  -13'd458,  
13'd1336,  13'd535,  13'd1555,  13'd949,  -13'd885,  13'd1029,  13'd27,  -13'd32,  13'd983,  -13'd603,  -13'd339,  13'd321,  13'd596,  -13'd41,  -13'd532,  -13'd479,  

13'd38,  -13'd465,  -13'd625,  13'd13,  -13'd345,  13'd112,  -13'd153,  -13'd63,  13'd442,  -13'd419,  13'd273,  -13'd54,  -13'd203,  -13'd150,  -13'd124,  -13'd222,  
-13'd644,  13'd548,  13'd62,  -13'd974,  13'd91,  -13'd611,  13'd263,  -13'd384,  13'd366,  13'd12,  13'd32,  -13'd508,  13'd121,  -13'd17,  -13'd408,  13'd201,  
13'd276,  13'd26,  -13'd79,  -13'd399,  13'd227,  -13'd565,  -13'd458,  -13'd69,  -13'd193,  -13'd77,  -13'd191,  -13'd451,  -13'd722,  -13'd109,  -13'd61,  -13'd508,  
13'd399,  -13'd431,  -13'd251,  -13'd511,  -13'd77,  -13'd236,  13'd123,  -13'd291,  -13'd577,  -13'd133,  -13'd742,  13'd132,  -13'd332,  -13'd757,  -13'd98,  13'd73,  
-13'd14,  -13'd521,  13'd31,  13'd573,  -13'd108,  13'd579,  -13'd848,  13'd567,  -13'd378,  13'd365,  13'd181,  -13'd118,  -13'd503,  13'd203,  -13'd52,  13'd125,  
13'd337,  -13'd443,  13'd358,  13'd445,  -13'd690,  13'd93,  13'd392,  -13'd411,  -13'd765,  -13'd439,  13'd222,  -13'd303,  -13'd262,  13'd271,  13'd41,  13'd254,  
-13'd117,  -13'd435,  -13'd77,  -13'd52,  -13'd689,  -13'd138,  -13'd171,  -13'd53,  -13'd124,  -13'd475,  -13'd245,  -13'd507,  13'd176,  13'd426,  13'd186,  -13'd350,  
-13'd775,  -13'd24,  -13'd366,  -13'd342,  -13'd400,  -13'd120,  -13'd301,  -13'd454,  -13'd523,  -13'd508,  -13'd295,  13'd379,  13'd138,  -13'd155,  -13'd842,  13'd297,  
-13'd326,  -13'd110,  -13'd187,  13'd99,  13'd397,  -13'd335,  -13'd146,  -13'd232,  -13'd529,  -13'd277,  13'd201,  13'd424,  -13'd94,  -13'd158,  13'd85,  -13'd241,  
13'd60,  -13'd432,  -13'd378,  -13'd459,  -13'd241,  -13'd142,  -13'd382,  13'd162,  13'd158,  -13'd339,  -13'd450,  13'd129,  13'd495,  13'd412,  13'd315,  -13'd228,  
-13'd747,  13'd73,  -13'd14,  -13'd382,  13'd176,  13'd94,  -13'd265,  -13'd153,  13'd140,  -13'd115,  -13'd428,  13'd90,  13'd164,  13'd189,  -13'd254,  -13'd690,  
-13'd175,  -13'd616,  13'd17,  -13'd824,  -13'd578,  13'd168,  13'd345,  -13'd230,  -13'd212,  13'd155,  13'd544,  -13'd18,  13'd270,  13'd159,  -13'd905,  -13'd781,  
13'd161,  -13'd773,  13'd640,  -13'd18,  -13'd546,  -13'd639,  13'd194,  -13'd51,  -13'd523,  13'd402,  -13'd239,  13'd290,  13'd19,  13'd593,  13'd30,  -13'd558,  
13'd699,  13'd86,  13'd22,  -13'd684,  -13'd427,  -13'd189,  -13'd146,  -13'd357,  -13'd45,  13'd301,  13'd331,  -13'd251,  -13'd106,  -13'd399,  13'd254,  13'd104,  
-13'd156,  -13'd5,  13'd124,  13'd408,  -13'd234,  -13'd421,  -13'd582,  -13'd331,  -13'd186,  -13'd34,  -13'd142,  13'd529,  13'd156,  -13'd184,  13'd238,  -13'd116,  
13'd650,  -13'd774,  -13'd461,  13'd192,  -13'd889,  13'd92,  13'd306,  -13'd591,  -13'd133,  -13'd476,  13'd361,  13'd156,  -13'd232,  -13'd382,  -13'd397,  -13'd122,  
13'd116,  13'd231,  13'd184,  13'd366,  -13'd209,  -13'd676,  13'd445,  13'd318,  -13'd209,  13'd120,  -13'd287,  13'd235,  13'd110,  -13'd558,  -13'd84,  -13'd393,  
-13'd288,  -13'd208,  -13'd153,  -13'd586,  -13'd169,  -13'd215,  13'd209,  -13'd134,  -13'd57,  -13'd125,  13'd522,  -13'd554,  -13'd109,  -13'd18,  -13'd423,  13'd233,  
-13'd575,  13'd429,  13'd550,  13'd40,  13'd195,  -13'd360,  -13'd679,  -13'd271,  -13'd478,  -13'd649,  13'd291,  -13'd373,  13'd31,  13'd94,  13'd492,  13'd150,  
-13'd417,  -13'd439,  -13'd501,  -13'd612,  -13'd317,  13'd309,  13'd440,  13'd3,  -13'd655,  13'd160,  13'd293,  13'd563,  -13'd235,  -13'd546,  13'd70,  -13'd124,  
13'd203,  -13'd544,  13'd218,  -13'd347,  -13'd402,  -13'd485,  13'd277,  13'd267,  -13'd127,  -13'd383,  -13'd73,  13'd426,  -13'd49,  -13'd198,  13'd153,  -13'd74,  
-13'd254,  -13'd869,  -13'd35,  13'd12,  -13'd118,  13'd282,  -13'd461,  -13'd776,  -13'd113,  -13'd141,  13'd314,  -13'd350,  13'd56,  13'd41,  -13'd728,  -13'd59,  
-13'd351,  -13'd230,  13'd506,  13'd195,  13'd488,  -13'd189,  -13'd536,  -13'd164,  13'd34,  -13'd223,  13'd599,  -13'd674,  -13'd620,  -13'd9,  13'd132,  -13'd690,  
-13'd233,  -13'd20,  13'd345,  -13'd87,  13'd375,  13'd195,  -13'd324,  13'd89,  -13'd90,  13'd5,  13'd199,  -13'd94,  -13'd537,  -13'd824,  -13'd14,  13'd99,  
-13'd557,  -13'd8,  -13'd165,  -13'd300,  13'd50,  -13'd693,  13'd420,  13'd202,  -13'd644,  13'd32,  -13'd4,  -13'd1023,  13'd137,  13'd171,  -13'd250,  13'd99,  

13'd172,  -13'd416,  13'd328,  -13'd842,  -13'd248,  -13'd357,  13'd730,  -13'd29,  13'd33,  -13'd93,  -13'd788,  -13'd100,  -13'd239,  13'd174,  -13'd121,  -13'd136,  
13'd886,  13'd583,  -13'd52,  -13'd758,  -13'd854,  13'd927,  13'd1071,  13'd193,  13'd133,  -13'd53,  -13'd92,  -13'd0,  13'd680,  13'd1045,  13'd47,  -13'd56,  
13'd141,  -13'd281,  -13'd212,  13'd158,  -13'd154,  13'd259,  13'd826,  -13'd27,  13'd129,  -13'd411,  13'd570,  13'd219,  13'd117,  13'd370,  13'd2,  13'd371,  
13'd475,  13'd492,  13'd217,  13'd136,  13'd975,  13'd1187,  -13'd436,  13'd222,  13'd991,  13'd138,  13'd109,  -13'd310,  13'd395,  -13'd184,  13'd489,  -13'd16,  
13'd343,  13'd98,  13'd47,  -13'd617,  13'd25,  -13'd95,  -13'd193,  13'd693,  -13'd713,  13'd67,  13'd632,  13'd196,  13'd937,  -13'd402,  13'd199,  -13'd174,  
-13'd92,  -13'd910,  13'd297,  -13'd562,  -13'd10,  13'd337,  13'd504,  -13'd22,  -13'd378,  -13'd6,  13'd483,  -13'd271,  -13'd716,  13'd0,  13'd80,  13'd46,  
-13'd105,  13'd106,  13'd500,  -13'd717,  13'd603,  13'd55,  13'd394,  13'd250,  -13'd156,  -13'd58,  13'd921,  13'd282,  13'd439,  13'd429,  -13'd248,  -13'd110,  
13'd228,  -13'd90,  13'd945,  -13'd46,  -13'd226,  13'd624,  13'd236,  13'd365,  13'd313,  -13'd165,  -13'd15,  -13'd851,  -13'd236,  -13'd92,  13'd229,  -13'd489,  
13'd526,  13'd549,  -13'd19,  -13'd378,  -13'd20,  13'd480,  -13'd934,  -13'd258,  13'd123,  -13'd123,  13'd291,  -13'd46,  13'd189,  -13'd501,  -13'd745,  13'd564,  
-13'd865,  -13'd484,  13'd1116,  13'd313,  -13'd408,  13'd79,  -13'd46,  -13'd367,  -13'd18,  13'd281,  13'd2,  13'd773,  -13'd153,  -13'd245,  13'd595,  13'd919,  
-13'd456,  13'd759,  -13'd141,  -13'd237,  -13'd916,  -13'd848,  13'd277,  13'd20,  -13'd1367,  -13'd431,  -13'd605,  13'd2,  -13'd520,  13'd167,  13'd544,  13'd210,  
13'd656,  -13'd655,  13'd88,  -13'd237,  -13'd504,  -13'd646,  -13'd408,  -13'd894,  -13'd378,  -13'd819,  -13'd2,  13'd399,  -13'd728,  13'd358,  -13'd3,  13'd46,  
-13'd156,  -13'd79,  -13'd20,  13'd52,  -13'd227,  -13'd424,  -13'd2,  13'd123,  13'd343,  -13'd484,  -13'd186,  -13'd222,  -13'd597,  -13'd416,  13'd354,  13'd7,  
-13'd1050,  13'd393,  -13'd328,  -13'd358,  13'd663,  -13'd373,  13'd567,  -13'd465,  -13'd294,  13'd325,  13'd65,  13'd196,  -13'd340,  -13'd197,  -13'd307,  -13'd390,  
-13'd485,  -13'd161,  13'd457,  -13'd151,  -13'd593,  13'd838,  13'd158,  -13'd41,  -13'd182,  13'd96,  -13'd63,  13'd267,  -13'd1816,  -13'd85,  -13'd204,  13'd31,  
13'd297,  13'd374,  13'd725,  -13'd527,  -13'd587,  -13'd204,  13'd351,  13'd174,  -13'd1050,  -13'd469,  -13'd873,  13'd43,  13'd3,  13'd645,  -13'd79,  13'd437,  
13'd522,  -13'd8,  13'd1111,  -13'd386,  -13'd203,  13'd673,  13'd967,  13'd589,  13'd111,  -13'd792,  -13'd504,  13'd206,  -13'd838,  13'd1014,  13'd488,  13'd65,  
13'd114,  -13'd26,  -13'd691,  13'd24,  -13'd54,  -13'd615,  13'd344,  13'd228,  -13'd811,  -13'd380,  -13'd158,  13'd105,  -13'd1174,  13'd164,  -13'd375,  -13'd435,  
-13'd798,  -13'd128,  -13'd509,  13'd236,  -13'd299,  -13'd224,  -13'd127,  -13'd361,  -13'd276,  -13'd215,  -13'd641,  13'd297,  13'd403,  13'd701,  13'd163,  -13'd338,  
-13'd101,  -13'd81,  -13'd164,  -13'd624,  13'd202,  13'd270,  13'd520,  -13'd315,  13'd1112,  13'd267,  -13'd261,  -13'd493,  -13'd811,  13'd278,  -13'd331,  -13'd1075,  
-13'd62,  -13'd525,  13'd264,  -13'd265,  -13'd132,  13'd27,  13'd92,  13'd229,  -13'd861,  13'd687,  -13'd583,  -13'd587,  -13'd123,  13'd1012,  -13'd136,  -13'd112,  
-13'd0,  -13'd406,  13'd189,  13'd830,  13'd438,  13'd944,  -13'd517,  13'd110,  -13'd228,  -13'd15,  -13'd93,  -13'd155,  -13'd286,  -13'd522,  13'd778,  13'd153,  
-13'd260,  13'd421,  -13'd553,  13'd585,  -13'd240,  -13'd86,  13'd205,  -13'd128,  13'd286,  13'd162,  -13'd88,  -13'd563,  13'd256,  13'd118,  13'd406,  -13'd752,  
-13'd538,  -13'd351,  -13'd14,  -13'd372,  13'd766,  -13'd886,  13'd132,  -13'd74,  13'd691,  13'd21,  13'd259,  13'd409,  -13'd8,  13'd60,  13'd56,  -13'd94,  
13'd365,  -13'd380,  -13'd470,  13'd561,  -13'd27,  13'd715,  -13'd287,  -13'd398,  13'd484,  13'd878,  -13'd748,  13'd775,  13'd309,  -13'd24,  13'd4,  -13'd221,  

-13'd1027,  13'd11,  -13'd348,  -13'd19,  13'd819,  13'd220,  -13'd260,  -13'd89,  13'd117,  -13'd513,  13'd130,  13'd329,  13'd678,  -13'd271,  13'd60,  13'd499,  
13'd7,  13'd369,  -13'd46,  -13'd26,  13'd1013,  -13'd371,  13'd217,  13'd18,  13'd609,  -13'd493,  -13'd452,  13'd532,  -13'd42,  13'd363,  -13'd15,  13'd197,  
-13'd84,  13'd825,  13'd63,  -13'd893,  13'd29,  -13'd3,  13'd188,  -13'd82,  -13'd678,  -13'd525,  -13'd601,  -13'd28,  -13'd372,  13'd1355,  -13'd8,  13'd466,  
-13'd510,  13'd611,  -13'd203,  13'd195,  13'd130,  13'd253,  13'd869,  -13'd24,  13'd205,  13'd159,  13'd61,  -13'd649,  -13'd299,  13'd1592,  13'd66,  13'd372,  
-13'd118,  13'd303,  -13'd254,  -13'd711,  13'd208,  13'd234,  13'd492,  13'd518,  13'd592,  13'd678,  13'd425,  -13'd302,  -13'd701,  13'd606,  13'd423,  -13'd596,  
-13'd328,  13'd118,  13'd248,  13'd12,  13'd183,  -13'd438,  13'd1220,  -13'd345,  -13'd293,  -13'd355,  13'd486,  13'd431,  13'd413,  -13'd163,  -13'd732,  13'd451,  
13'd149,  13'd72,  -13'd224,  -13'd63,  13'd131,  -13'd12,  13'd155,  -13'd53,  -13'd164,  13'd552,  -13'd123,  13'd342,  -13'd349,  -13'd103,  -13'd220,  -13'd222,  
13'd133,  -13'd492,  -13'd78,  -13'd802,  -13'd242,  -13'd389,  13'd122,  -13'd244,  -13'd218,  13'd480,  -13'd695,  13'd386,  -13'd377,  -13'd372,  -13'd296,  -13'd800,  
-13'd332,  -13'd689,  13'd910,  13'd428,  -13'd153,  13'd347,  13'd414,  -13'd912,  -13'd429,  13'd299,  13'd712,  13'd110,  13'd178,  13'd0,  -13'd114,  -13'd400,  
13'd431,  13'd727,  13'd323,  13'd177,  -13'd672,  13'd193,  13'd50,  -13'd264,  13'd362,  13'd256,  -13'd10,  13'd208,  13'd243,  -13'd756,  13'd54,  -13'd126,  
13'd475,  13'd435,  13'd108,  -13'd750,  -13'd776,  13'd84,  13'd255,  -13'd398,  -13'd331,  13'd340,  13'd909,  13'd428,  -13'd552,  -13'd273,  -13'd498,  13'd1,  
-13'd181,  13'd463,  -13'd467,  13'd663,  13'd259,  13'd817,  -13'd125,  13'd108,  13'd485,  -13'd536,  -13'd220,  13'd517,  13'd121,  -13'd94,  13'd515,  13'd758,  
-13'd53,  13'd330,  13'd333,  -13'd133,  -13'd252,  13'd155,  13'd20,  -13'd102,  13'd383,  13'd600,  13'd65,  -13'd123,  13'd368,  13'd441,  -13'd96,  13'd110,  
-13'd313,  13'd14,  13'd457,  13'd397,  -13'd496,  -13'd200,  -13'd223,  -13'd852,  13'd34,  13'd312,  13'd123,  13'd59,  13'd230,  13'd223,  -13'd145,  13'd727,  
13'd614,  -13'd421,  13'd120,  13'd642,  -13'd155,  13'd465,  13'd412,  -13'd201,  13'd212,  13'd329,  13'd543,  13'd370,  13'd165,  -13'd357,  -13'd719,  -13'd503,  
13'd616,  13'd462,  -13'd89,  -13'd294,  -13'd1037,  13'd350,  13'd372,  -13'd188,  -13'd714,  -13'd752,  13'd72,  13'd1035,  13'd558,  13'd291,  13'd324,  13'd812,  
13'd1149,  -13'd650,  13'd149,  13'd79,  13'd249,  13'd181,  13'd76,  -13'd74,  13'd420,  13'd340,  13'd101,  13'd163,  -13'd437,  13'd245,  13'd824,  -13'd460,  
13'd264,  13'd93,  -13'd587,  13'd523,  13'd337,  -13'd139,  -13'd203,  13'd330,  13'd225,  13'd182,  13'd13,  13'd499,  13'd789,  -13'd532,  -13'd422,  13'd596,  
13'd217,  13'd242,  -13'd133,  -13'd223,  13'd595,  -13'd668,  -13'd876,  -13'd366,  13'd117,  13'd38,  13'd156,  -13'd609,  13'd279,  -13'd435,  13'd218,  13'd220,  
13'd460,  13'd500,  13'd266,  -13'd184,  13'd218,  13'd42,  -13'd202,  13'd242,  13'd264,  -13'd151,  13'd678,  13'd389,  13'd6,  13'd299,  -13'd410,  13'd672,  
13'd838,  13'd0,  13'd228,  13'd898,  13'd392,  13'd176,  -13'd29,  13'd478,  -13'd350,  13'd840,  -13'd118,  13'd217,  13'd407,  13'd688,  13'd32,  13'd458,  
13'd193,  -13'd193,  13'd294,  -13'd86,  13'd425,  13'd480,  -13'd577,  13'd759,  -13'd1267,  -13'd247,  13'd604,  -13'd448,  13'd194,  13'd483,  -13'd465,  13'd22,  
13'd280,  -13'd118,  -13'd241,  13'd254,  -13'd481,  13'd728,  13'd369,  13'd639,  -13'd1068,  -13'd156,  -13'd139,  -13'd169,  13'd179,  -13'd966,  13'd281,  13'd377,  
13'd182,  -13'd71,  -13'd289,  -13'd152,  13'd607,  -13'd641,  -13'd162,  13'd273,  -13'd217,  13'd60,  -13'd222,  -13'd602,  13'd667,  -13'd9,  13'd368,  -13'd387,  
13'd151,  -13'd438,  -13'd982,  -13'd36,  13'd495,  13'd412,  13'd311,  13'd324,  -13'd468,  -13'd153,  13'd250,  13'd649,  13'd834,  -13'd366,  -13'd440,  13'd148,  

13'd1058,  13'd278,  13'd655,  13'd760,  -13'd226,  13'd474,  13'd1155,  13'd778,  -13'd45,  -13'd461,  13'd180,  -13'd285,  13'd159,  13'd1080,  -13'd100,  -13'd400,  
-13'd12,  13'd346,  13'd232,  13'd819,  -13'd528,  13'd379,  -13'd141,  -13'd66,  13'd374,  -13'd209,  13'd532,  13'd1047,  13'd56,  13'd444,  13'd43,  13'd523,  
-13'd382,  13'd140,  13'd221,  13'd293,  13'd572,  -13'd230,  13'd515,  -13'd54,  13'd708,  13'd1082,  13'd804,  13'd123,  13'd281,  13'd486,  -13'd468,  -13'd149,  
-13'd544,  -13'd400,  13'd1314,  13'd34,  -13'd405,  -13'd157,  -13'd719,  13'd683,  -13'd104,  13'd652,  -13'd319,  13'd527,  13'd263,  13'd704,  13'd617,  13'd68,  
-13'd428,  -13'd1385,  -13'd406,  -13'd324,  -13'd91,  -13'd659,  -13'd628,  -13'd391,  -13'd1300,  13'd200,  13'd228,  -13'd151,  -13'd3,  -13'd186,  -13'd455,  -13'd478,  
13'd252,  -13'd178,  13'd722,  13'd485,  -13'd779,  -13'd53,  -13'd403,  -13'd145,  13'd158,  13'd567,  -13'd147,  13'd134,  13'd496,  13'd66,  13'd114,  13'd353,  
-13'd273,  -13'd93,  13'd803,  13'd821,  -13'd565,  13'd351,  13'd301,  13'd458,  -13'd488,  13'd521,  13'd303,  -13'd705,  13'd583,  -13'd287,  13'd59,  13'd210,  
-13'd14,  13'd58,  -13'd684,  13'd610,  -13'd73,  13'd120,  -13'd631,  13'd194,  -13'd637,  -13'd558,  -13'd193,  -13'd289,  13'd896,  13'd217,  13'd602,  13'd306,  
-13'd494,  13'd330,  13'd358,  13'd471,  -13'd1025,  13'd159,  -13'd432,  13'd128,  -13'd690,  -13'd211,  -13'd497,  13'd39,  -13'd978,  13'd830,  13'd142,  -13'd364,  
-13'd183,  -13'd883,  13'd571,  -13'd79,  -13'd979,  -13'd29,  -13'd814,  13'd391,  -13'd311,  13'd278,  13'd363,  13'd362,  -13'd1016,  13'd710,  -13'd171,  -13'd984,  
13'd350,  13'd44,  -13'd643,  -13'd433,  13'd161,  13'd66,  13'd511,  -13'd75,  -13'd605,  -13'd98,  13'd1191,  -13'd654,  13'd370,  13'd165,  13'd151,  -13'd478,  
-13'd467,  13'd324,  -13'd618,  -13'd190,  -13'd657,  -13'd328,  -13'd1201,  -13'd137,  13'd125,  13'd149,  -13'd363,  -13'd830,  13'd303,  -13'd91,  13'd460,  -13'd235,  
-13'd602,  13'd516,  -13'd592,  13'd169,  13'd347,  -13'd759,  13'd266,  -13'd613,  13'd231,  -13'd507,  -13'd396,  -13'd243,  -13'd339,  13'd456,  -13'd220,  -13'd208,  
-13'd842,  13'd276,  13'd490,  -13'd277,  -13'd1056,  -13'd440,  -13'd221,  -13'd86,  -13'd696,  -13'd443,  13'd1202,  13'd290,  -13'd688,  -13'd235,  -13'd291,  -13'd350,  
13'd525,  13'd253,  13'd165,  -13'd77,  13'd208,  -13'd48,  -13'd348,  -13'd690,  -13'd561,  -13'd920,  -13'd114,  -13'd111,  -13'd393,  -13'd497,  13'd41,  -13'd167,  
-13'd69,  13'd66,  -13'd18,  -13'd636,  -13'd439,  -13'd676,  13'd362,  -13'd229,  13'd97,  -13'd89,  13'd24,  13'd49,  13'd225,  -13'd187,  -13'd116,  -13'd135,  
-13'd716,  -13'd317,  13'd602,  13'd135,  -13'd24,  -13'd529,  -13'd102,  -13'd467,  13'd259,  13'd285,  13'd312,  13'd1060,  -13'd420,  -13'd378,  13'd447,  13'd507,  
13'd58,  13'd108,  13'd727,  13'd170,  13'd413,  13'd698,  13'd631,  -13'd35,  13'd1270,  13'd1223,  -13'd954,  -13'd83,  -13'd199,  13'd736,  13'd299,  -13'd1020,  
13'd219,  13'd43,  13'd642,  13'd177,  -13'd299,  13'd173,  13'd146,  13'd16,  13'd217,  13'd110,  -13'd591,  13'd266,  -13'd530,  13'd314,  13'd474,  -13'd1088,  
13'd722,  -13'd563,  -13'd47,  -13'd63,  -13'd134,  -13'd206,  -13'd578,  -13'd340,  13'd328,  13'd510,  -13'd422,  13'd42,  13'd594,  -13'd179,  13'd368,  -13'd271,  
13'd410,  -13'd151,  13'd56,  13'd701,  -13'd400,  13'd86,  13'd882,  13'd449,  -13'd43,  -13'd654,  -13'd61,  13'd10,  -13'd35,  -13'd390,  -13'd8,  -13'd83,  
-13'd507,  -13'd120,  13'd254,  13'd1025,  -13'd406,  13'd1057,  13'd134,  -13'd137,  13'd875,  -13'd63,  13'd142,  13'd521,  13'd351,  13'd318,  -13'd440,  13'd103,  
13'd337,  -13'd136,  13'd85,  13'd888,  13'd975,  13'd677,  13'd305,  -13'd163,  -13'd440,  13'd214,  13'd627,  -13'd424,  13'd632,  13'd249,  -13'd27,  13'd162,  
-13'd651,  13'd497,  -13'd962,  13'd667,  13'd180,  13'd133,  -13'd514,  -13'd20,  13'd264,  13'd458,  13'd272,  -13'd305,  13'd457,  -13'd741,  13'd510,  13'd99,  
-13'd741,  -13'd678,  13'd140,  13'd621,  13'd128,  13'd9,  -13'd213,  -13'd247,  -13'd212,  13'd1109,  13'd679,  13'd253,  13'd426,  -13'd1127,  13'd430,  -13'd154,  

-13'd494,  13'd66,  13'd401,  13'd652,  -13'd466,  -13'd95,  -13'd476,  13'd294,  -13'd279,  13'd284,  -13'd263,  -13'd877,  13'd948,  -13'd315,  13'd627,  13'd107,  
13'd33,  -13'd145,  13'd104,  13'd87,  13'd164,  -13'd643,  -13'd539,  -13'd0,  13'd486,  -13'd13,  13'd24,  13'd638,  -13'd282,  -13'd121,  13'd264,  -13'd45,  
13'd85,  -13'd140,  13'd578,  13'd168,  13'd143,  -13'd307,  -13'd91,  13'd146,  -13'd185,  13'd110,  13'd140,  13'd98,  13'd646,  13'd662,  -13'd203,  -13'd661,  
-13'd17,  13'd26,  -13'd378,  -13'd399,  13'd45,  -13'd294,  13'd33,  -13'd336,  -13'd32,  -13'd348,  -13'd301,  13'd107,  -13'd293,  13'd75,  -13'd214,  -13'd562,  
13'd643,  13'd367,  -13'd192,  13'd45,  -13'd305,  13'd58,  -13'd257,  -13'd269,  -13'd555,  -13'd273,  13'd112,  13'd686,  -13'd478,  13'd48,  -13'd105,  -13'd193,  
-13'd36,  13'd360,  13'd2,  13'd219,  13'd355,  13'd650,  -13'd641,  -13'd305,  13'd133,  13'd145,  -13'd116,  13'd686,  -13'd192,  -13'd292,  13'd365,  -13'd324,  
-13'd206,  -13'd163,  13'd291,  13'd235,  13'd670,  -13'd399,  13'd36,  13'd184,  13'd286,  -13'd323,  -13'd339,  13'd404,  13'd590,  -13'd251,  13'd124,  -13'd154,  
-13'd388,  13'd242,  -13'd404,  13'd637,  -13'd76,  -13'd197,  13'd342,  -13'd787,  13'd193,  -13'd154,  13'd202,  -13'd0,  13'd498,  13'd655,  -13'd119,  13'd289,  
-13'd193,  -13'd210,  -13'd56,  -13'd89,  13'd906,  13'd69,  13'd143,  -13'd61,  13'd938,  -13'd226,  13'd151,  -13'd170,  13'd25,  -13'd155,  -13'd85,  -13'd629,  
13'd1422,  13'd163,  -13'd604,  13'd753,  13'd659,  13'd265,  -13'd93,  13'd121,  -13'd33,  13'd676,  -13'd78,  13'd134,  13'd933,  13'd311,  13'd125,  13'd44,  
-13'd567,  13'd244,  -13'd136,  13'd282,  13'd260,  13'd690,  -13'd321,  13'd306,  13'd48,  -13'd485,  13'd46,  -13'd397,  -13'd147,  13'd67,  13'd498,  13'd480,  
-13'd139,  -13'd74,  -13'd24,  13'd203,  13'd106,  -13'd257,  -13'd247,  13'd828,  -13'd662,  13'd322,  -13'd460,  13'd697,  13'd529,  -13'd834,  13'd360,  13'd602,  
-13'd656,  13'd305,  -13'd385,  13'd379,  -13'd429,  13'd371,  13'd784,  -13'd242,  13'd182,  -13'd240,  13'd834,  -13'd161,  13'd1087,  13'd59,  -13'd453,  -13'd94,  
-13'd216,  -13'd509,  -13'd351,  13'd823,  -13'd192,  13'd520,  -13'd85,  -13'd112,  13'd605,  -13'd10,  13'd725,  -13'd0,  13'd655,  -13'd300,  -13'd148,  13'd325,  
-13'd935,  -13'd138,  13'd8,  13'd178,  -13'd84,  13'd279,  -13'd807,  13'd356,  13'd283,  -13'd350,  13'd172,  -13'd505,  13'd607,  13'd192,  13'd458,  -13'd302,  
-13'd330,  13'd549,  -13'd335,  -13'd446,  13'd654,  -13'd620,  -13'd890,  -13'd373,  -13'd97,  13'd1019,  13'd619,  -13'd544,  -13'd400,  13'd309,  -13'd891,  -13'd293,  
13'd101,  13'd830,  -13'd327,  -13'd224,  -13'd169,  13'd321,  -13'd353,  13'd244,  13'd110,  13'd411,  13'd485,  -13'd630,  13'd378,  -13'd1596,  -13'd631,  -13'd202,  
-13'd129,  13'd389,  -13'd858,  -13'd665,  13'd393,  -13'd178,  13'd88,  -13'd448,  13'd328,  -13'd101,  13'd161,  -13'd703,  -13'd209,  -13'd569,  -13'd380,  13'd755,  
-13'd669,  13'd661,  -13'd135,  -13'd427,  13'd924,  -13'd328,  13'd750,  -13'd465,  13'd937,  13'd290,  -13'd9,  13'd531,  -13'd85,  -13'd334,  13'd525,  13'd624,  
-13'd515,  13'd229,  -13'd985,  13'd133,  13'd28,  -13'd70,  13'd357,  13'd578,  -13'd150,  -13'd530,  13'd11,  13'd157,  -13'd527,  -13'd414,  -13'd592,  -13'd351,  
13'd259,  13'd59,  -13'd1116,  13'd228,  -13'd78,  -13'd332,  13'd1062,  -13'd810,  13'd504,  13'd219,  13'd316,  13'd640,  13'd157,  -13'd239,  -13'd488,  13'd170,  
13'd97,  13'd408,  -13'd550,  -13'd833,  13'd829,  -13'd457,  13'd378,  -13'd564,  13'd397,  13'd384,  -13'd67,  13'd218,  -13'd161,  -13'd648,  -13'd919,  -13'd41,  
13'd503,  13'd840,  13'd131,  -13'd1221,  13'd1172,  -13'd205,  13'd383,  -13'd616,  -13'd62,  13'd1537,  -13'd821,  -13'd90,  -13'd818,  13'd711,  -13'd599,  13'd314,  
-13'd513,  13'd175,  13'd275,  13'd10,  13'd363,  -13'd308,  13'd943,  -13'd669,  13'd86,  -13'd676,  -13'd928,  -13'd161,  -13'd106,  13'd459,  13'd10,  -13'd497,  
13'd33,  -13'd80,  13'd887,  -13'd381,  -13'd433,  13'd271,  13'd270,  -13'd511,  13'd677,  13'd355,  -13'd654,  13'd183,  -13'd497,  13'd329,  13'd34,  -13'd104,  

-13'd1343,  -13'd442,  -13'd679,  13'd297,  13'd154,  13'd48,  -13'd800,  13'd337,  13'd317,  -13'd58,  -13'd503,  -13'd224,  13'd202,  -13'd390,  -13'd157,  13'd485,  
13'd165,  -13'd622,  13'd660,  -13'd502,  13'd202,  -13'd433,  13'd25,  13'd202,  -13'd15,  -13'd610,  -13'd676,  -13'd643,  -13'd52,  13'd415,  -13'd434,  -13'd35,  
-13'd708,  -13'd311,  13'd65,  13'd197,  -13'd325,  -13'd448,  -13'd21,  -13'd80,  -13'd690,  13'd44,  -13'd320,  -13'd398,  -13'd191,  13'd1622,  13'd97,  -13'd1011,  
13'd402,  -13'd523,  13'd784,  -13'd124,  -13'd604,  -13'd225,  -13'd48,  13'd179,  13'd34,  -13'd505,  13'd145,  -13'd63,  -13'd866,  -13'd36,  13'd217,  -13'd1053,  
13'd743,  -13'd4,  -13'd220,  13'd703,  -13'd404,  13'd699,  -13'd408,  13'd272,  13'd321,  13'd389,  13'd163,  13'd13,  13'd698,  -13'd573,  13'd323,  13'd620,  
-13'd261,  13'd381,  -13'd238,  13'd530,  13'd426,  -13'd261,  -13'd780,  -13'd605,  -13'd558,  13'd192,  -13'd119,  13'd135,  -13'd291,  13'd218,  13'd8,  -13'd186,  
13'd40,  -13'd532,  -13'd10,  -13'd506,  13'd473,  -13'd111,  13'd147,  13'd110,  -13'd138,  13'd232,  -13'd214,  13'd610,  -13'd982,  13'd274,  13'd165,  13'd22,  
13'd346,  13'd657,  13'd708,  13'd373,  13'd30,  13'd229,  -13'd649,  13'd428,  13'd294,  13'd219,  13'd40,  -13'd242,  -13'd21,  13'd940,  13'd257,  -13'd477,  
13'd7,  13'd108,  -13'd133,  13'd467,  -13'd578,  13'd629,  -13'd603,  13'd792,  -13'd517,  -13'd169,  -13'd5,  -13'd573,  13'd482,  -13'd44,  13'd46,  -13'd535,  
13'd760,  13'd263,  -13'd383,  13'd320,  13'd8,  13'd381,  -13'd669,  -13'd242,  -13'd254,  13'd1173,  13'd361,  -13'd496,  13'd716,  -13'd579,  13'd389,  13'd618,  
13'd91,  -13'd241,  13'd95,  13'd400,  -13'd897,  13'd538,  -13'd1041,  13'd438,  13'd404,  13'd13,  13'd686,  13'd398,  13'd265,  -13'd183,  13'd106,  -13'd71,  
13'd245,  -13'd886,  13'd141,  13'd285,  13'd579,  13'd177,  13'd23,  13'd209,  13'd715,  13'd34,  13'd477,  13'd557,  13'd343,  -13'd260,  13'd446,  13'd63,  
-13'd347,  13'd295,  13'd830,  13'd100,  -13'd336,  -13'd425,  13'd110,  -13'd224,  13'd519,  13'd73,  13'd264,  13'd883,  13'd36,  13'd905,  13'd110,  -13'd238,  
-13'd798,  -13'd30,  13'd577,  13'd115,  -13'd200,  13'd0,  13'd543,  -13'd61,  -13'd295,  13'd633,  13'd737,  13'd151,  -13'd124,  -13'd282,  13'd104,  -13'd785,  
-13'd839,  -13'd450,  13'd131,  13'd864,  13'd89,  13'd40,  -13'd691,  -13'd401,  13'd4,  13'd200,  13'd26,  -13'd85,  -13'd250,  -13'd439,  13'd204,  -13'd145,  
13'd443,  13'd266,  13'd204,  -13'd108,  -13'd96,  13'd131,  13'd514,  13'd201,  13'd498,  13'd228,  13'd1528,  -13'd573,  13'd903,  -13'd104,  13'd120,  -13'd33,  
-13'd277,  13'd307,  13'd22,  13'd513,  -13'd344,  13'd313,  13'd628,  13'd494,  -13'd45,  13'd158,  13'd7,  13'd493,  -13'd66,  -13'd103,  13'd103,  -13'd493,  
13'd145,  -13'd176,  13'd62,  -13'd188,  -13'd240,  13'd220,  -13'd571,  13'd6,  13'd653,  -13'd239,  13'd398,  -13'd443,  13'd360,  13'd1426,  13'd174,  -13'd74,  
-13'd594,  -13'd217,  13'd431,  -13'd46,  13'd179,  -13'd628,  13'd81,  13'd239,  13'd141,  -13'd372,  13'd390,  -13'd331,  13'd187,  13'd175,  13'd483,  13'd563,  
13'd418,  13'd595,  13'd1258,  13'd247,  -13'd324,  13'd520,  -13'd0,  -13'd3,  -13'd1,  13'd57,  13'd127,  13'd1035,  -13'd79,  -13'd35,  13'd125,  13'd215,  
13'd41,  13'd268,  -13'd619,  -13'd318,  -13'd393,  -13'd502,  13'd1554,  -13'd456,  13'd337,  -13'd838,  13'd494,  -13'd302,  -13'd130,  -13'd116,  13'd103,  13'd429,  
13'd370,  13'd75,  13'd147,  -13'd272,  13'd186,  13'd382,  13'd882,  13'd18,  13'd355,  13'd402,  -13'd119,  13'd385,  -13'd180,  13'd460,  -13'd268,  -13'd448,  
-13'd29,  -13'd205,  -13'd542,  -13'd592,  13'd344,  13'd25,  -13'd250,  13'd302,  -13'd93,  -13'd548,  13'd218,  13'd57,  -13'd425,  13'd909,  -13'd249,  13'd652,  
-13'd1318,  -13'd107,  13'd375,  -13'd127,  -13'd321,  13'd20,  13'd269,  13'd428,  13'd345,  13'd84,  -13'd743,  13'd518,  -13'd117,  13'd48,  13'd807,  13'd315,  
13'd1310,  13'd1022,  13'd818,  -13'd658,  13'd54,  13'd111,  -13'd532,  -13'd172,  -13'd314,  -13'd56,  13'd667,  13'd222,  13'd241,  -13'd197,  -13'd177,  13'd620,  

13'd3,  13'd566,  -13'd734,  13'd444,  -13'd422,  13'd598,  -13'd831,  -13'd323,  -13'd9,  13'd380,  13'd869,  13'd133,  13'd921,  -13'd394,  -13'd45,  -13'd503,  
13'd236,  -13'd283,  13'd9,  13'd246,  13'd205,  13'd727,  -13'd299,  -13'd735,  13'd311,  13'd113,  -13'd141,  13'd253,  13'd580,  -13'd970,  -13'd508,  -13'd106,  
13'd511,  -13'd291,  -13'd337,  -13'd170,  13'd628,  13'd664,  13'd323,  -13'd598,  -13'd607,  -13'd400,  13'd414,  13'd100,  13'd646,  -13'd261,  -13'd763,  -13'd520,  
13'd506,  13'd904,  13'd223,  13'd434,  13'd576,  13'd282,  -13'd250,  13'd161,  13'd489,  -13'd97,  13'd314,  -13'd173,  -13'd659,  13'd697,  13'd307,  13'd383,  
-13'd207,  13'd160,  13'd420,  13'd55,  -13'd766,  -13'd60,  -13'd212,  -13'd182,  -13'd139,  -13'd4,  -13'd364,  -13'd397,  -13'd1363,  -13'd931,  13'd679,  -13'd357,  
13'd226,  13'd285,  -13'd1213,  13'd59,  -13'd380,  13'd51,  13'd340,  13'd249,  13'd475,  -13'd367,  13'd790,  13'd259,  13'd376,  -13'd612,  -13'd712,  -13'd39,  
13'd103,  13'd294,  -13'd543,  13'd286,  -13'd470,  -13'd252,  13'd234,  13'd307,  -13'd138,  13'd21,  13'd520,  13'd581,  13'd836,  -13'd736,  -13'd1133,  13'd335,  
13'd591,  13'd856,  -13'd202,  -13'd503,  -13'd56,  -13'd147,  13'd594,  -13'd867,  13'd398,  -13'd546,  13'd163,  13'd163,  13'd449,  13'd819,  -13'd249,  13'd918,  
-13'd57,  13'd732,  13'd638,  -13'd843,  13'd562,  13'd405,  13'd250,  13'd110,  -13'd113,  13'd124,  -13'd241,  -13'd415,  -13'd135,  13'd1082,  -13'd533,  -13'd346,  
13'd164,  13'd470,  13'd477,  13'd246,  -13'd594,  13'd151,  13'd575,  13'd587,  -13'd473,  -13'd7,  13'd210,  -13'd377,  -13'd1052,  -13'd119,  13'd63,  -13'd1121,  
-13'd309,  -13'd706,  -13'd474,  -13'd943,  -13'd173,  -13'd948,  13'd464,  -13'd217,  -13'd270,  -13'd258,  13'd664,  -13'd292,  -13'd586,  -13'd361,  13'd403,  -13'd434,  
-13'd163,  -13'd833,  -13'd458,  13'd160,  -13'd791,  -13'd163,  -13'd603,  -13'd637,  13'd157,  13'd10,  13'd421,  13'd36,  -13'd375,  13'd178,  -13'd1232,  13'd449,  
-13'd5,  -13'd180,  -13'd704,  -13'd862,  13'd706,  -13'd492,  13'd356,  -13'd490,  13'd369,  13'd873,  13'd64,  -13'd323,  13'd254,  13'd445,  -13'd338,  -13'd344,  
13'd60,  13'd287,  13'd484,  -13'd838,  13'd261,  -13'd418,  13'd291,  -13'd647,  13'd407,  13'd62,  13'd112,  -13'd162,  13'd16,  13'd1046,  -13'd516,  -13'd291,  
13'd1230,  13'd602,  -13'd50,  13'd357,  -13'd361,  -13'd11,  13'd572,  13'd325,  13'd470,  13'd246,  13'd549,  -13'd343,  -13'd162,  -13'd506,  -13'd65,  -13'd194,  
-13'd345,  -13'd222,  13'd168,  13'd356,  -13'd488,  -13'd223,  -13'd86,  -13'd583,  -13'd76,  -13'd333,  -13'd118,  13'd216,  -13'd577,  -13'd208,  -13'd20,  -13'd645,  
13'd212,  -13'd877,  -13'd583,  -13'd693,  13'd332,  -13'd501,  -13'd585,  -13'd630,  13'd501,  -13'd360,  13'd232,  13'd364,  13'd121,  -13'd195,  -13'd511,  -13'd599,  
-13'd36,  -13'd540,  13'd60,  -13'd300,  13'd147,  -13'd962,  13'd240,  -13'd508,  13'd611,  13'd138,  -13'd492,  13'd760,  -13'd443,  -13'd341,  -13'd245,  -13'd346,  
13'd180,  -13'd503,  13'd228,  -13'd19,  13'd224,  -13'd102,  -13'd417,  13'd117,  13'd837,  13'd147,  -13'd592,  -13'd488,  13'd153,  13'd902,  13'd39,  -13'd654,  
13'd67,  -13'd133,  -13'd1013,  -13'd473,  -13'd221,  13'd636,  -13'd95,  13'd531,  13'd1212,  13'd545,  13'd169,  13'd388,  13'd369,  -13'd969,  13'd817,  -13'd454,  
13'd507,  13'd0,  13'd397,  13'd423,  -13'd991,  13'd207,  -13'd108,  -13'd156,  13'd24,  -13'd995,  13'd317,  13'd105,  13'd261,  -13'd182,  -13'd54,  13'd47,  
13'd249,  -13'd682,  -13'd743,  13'd742,  -13'd747,  13'd456,  -13'd218,  13'd195,  13'd32,  -13'd53,  13'd676,  13'd9,  13'd182,  -13'd49,  -13'd138,  13'd666,  
13'd394,  13'd181,  13'd9,  13'd468,  -13'd577,  13'd792,  13'd82,  13'd185,  13'd155,  -13'd376,  13'd819,  -13'd144,  13'd867,  13'd130,  13'd401,  -13'd39,  
-13'd717,  13'd242,  13'd448,  13'd341,  13'd766,  13'd536,  -13'd520,  -13'd143,  -13'd93,  13'd1001,  13'd285,  -13'd201,  13'd302,  -13'd961,  13'd295,  13'd532,  
-13'd667,  -13'd389,  13'd250,  13'd293,  -13'd60,  13'd656,  13'd99,  13'd257,  13'd294,  13'd816,  13'd748,  13'd640,  13'd392,  -13'd246,  13'd160,  13'd306,  

-13'd541,  -13'd555,  13'd140,  13'd436,  -13'd50,  13'd168,  -13'd110,  -13'd468,  13'd138,  13'd151,  13'd138,  -13'd61,  -13'd595,  -13'd234,  13'd559,  13'd97,  
13'd64,  13'd218,  13'd204,  -13'd276,  13'd144,  -13'd600,  13'd196,  -13'd275,  -13'd231,  -13'd261,  -13'd4,  -13'd660,  13'd195,  13'd333,  -13'd15,  -13'd376,  
13'd396,  -13'd216,  -13'd568,  13'd157,  13'd337,  -13'd866,  -13'd23,  13'd18,  -13'd70,  -13'd205,  -13'd209,  13'd137,  13'd318,  13'd559,  13'd92,  -13'd280,  
13'd389,  -13'd165,  -13'd273,  13'd385,  -13'd487,  13'd519,  -13'd430,  13'd45,  -13'd146,  13'd218,  -13'd348,  -13'd239,  -13'd509,  13'd528,  13'd291,  -13'd539,  
13'd479,  13'd21,  13'd63,  -13'd403,  -13'd46,  -13'd111,  13'd15,  13'd741,  13'd244,  -13'd580,  -13'd368,  13'd189,  13'd3,  13'd301,  -13'd111,  -13'd633,  
13'd17,  -13'd40,  13'd639,  -13'd507,  -13'd364,  13'd735,  -13'd31,  -13'd228,  -13'd279,  13'd514,  -13'd427,  13'd285,  13'd177,  -13'd583,  -13'd219,  -13'd136,  
13'd369,  13'd409,  -13'd125,  -13'd214,  -13'd125,  -13'd488,  -13'd390,  -13'd286,  13'd671,  -13'd674,  -13'd239,  -13'd513,  -13'd364,  -13'd879,  13'd615,  -13'd835,  
13'd131,  13'd156,  -13'd105,  -13'd396,  -13'd386,  -13'd205,  -13'd130,  13'd9,  -13'd105,  -13'd477,  13'd455,  13'd386,  13'd396,  -13'd123,  13'd213,  13'd290,  
13'd324,  13'd483,  13'd187,  -13'd285,  -13'd75,  13'd54,  -13'd756,  13'd405,  -13'd419,  -13'd423,  13'd206,  -13'd853,  13'd208,  -13'd185,  -13'd366,  -13'd838,  
-13'd128,  -13'd151,  13'd102,  13'd134,  -13'd377,  13'd142,  -13'd93,  -13'd59,  -13'd560,  -13'd324,  -13'd450,  13'd494,  13'd153,  -13'd311,  13'd290,  -13'd562,  
13'd386,  13'd136,  13'd209,  13'd231,  13'd148,  13'd149,  -13'd297,  13'd4,  -13'd106,  -13'd298,  -13'd120,  13'd43,  13'd111,  -13'd390,  -13'd192,  13'd31,  
13'd383,  -13'd287,  13'd385,  13'd739,  -13'd290,  13'd56,  -13'd649,  -13'd628,  13'd139,  -13'd121,  -13'd175,  -13'd609,  13'd695,  -13'd27,  -13'd145,  -13'd226,  
13'd217,  13'd178,  -13'd343,  -13'd395,  13'd90,  -13'd737,  13'd382,  -13'd581,  13'd544,  13'd565,  13'd423,  -13'd387,  -13'd155,  -13'd278,  -13'd759,  -13'd168,  
13'd102,  -13'd474,  13'd204,  13'd465,  -13'd307,  -13'd228,  -13'd80,  13'd264,  13'd634,  -13'd381,  13'd138,  -13'd463,  13'd219,  13'd379,  13'd686,  13'd273,  
13'd330,  -13'd629,  13'd84,  13'd126,  -13'd229,  13'd26,  13'd397,  13'd267,  -13'd154,  -13'd318,  -13'd108,  -13'd177,  -13'd414,  13'd333,  13'd54,  -13'd285,  
-13'd149,  13'd50,  13'd572,  -13'd243,  -13'd279,  -13'd481,  13'd108,  -13'd20,  13'd40,  13'd202,  -13'd210,  -13'd256,  -13'd265,  -13'd274,  -13'd48,  -13'd282,  
13'd248,  -13'd148,  -13'd329,  -13'd536,  13'd179,  -13'd501,  -13'd135,  13'd160,  -13'd384,  13'd277,  -13'd210,  13'd202,  -13'd603,  13'd438,  -13'd143,  -13'd117,  
-13'd94,  -13'd341,  -13'd58,  -13'd56,  -13'd20,  13'd106,  -13'd416,  -13'd467,  13'd90,  -13'd382,  -13'd16,  -13'd465,  13'd1,  -13'd111,  -13'd489,  13'd155,  
13'd250,  -13'd139,  -13'd290,  -13'd363,  -13'd629,  13'd397,  -13'd4,  -13'd226,  -13'd78,  13'd35,  13'd152,  -13'd588,  -13'd160,  -13'd888,  -13'd82,  -13'd112,  
13'd774,  -13'd468,  -13'd271,  -13'd258,  -13'd261,  -13'd56,  -13'd57,  -13'd140,  13'd248,  -13'd36,  13'd29,  13'd86,  13'd522,  13'd374,  -13'd31,  -13'd822,  
13'd177,  -13'd45,  -13'd76,  -13'd708,  -13'd194,  13'd630,  -13'd45,  -13'd114,  -13'd10,  13'd561,  -13'd610,  -13'd130,  -13'd432,  13'd261,  13'd334,  -13'd185,  
-13'd138,  -13'd871,  -13'd517,  -13'd44,  -13'd329,  -13'd215,  -13'd221,  13'd442,  13'd328,  -13'd18,  -13'd509,  -13'd356,  -13'd660,  -13'd742,  -13'd3,  13'd456,  
-13'd240,  -13'd145,  13'd294,  13'd59,  13'd152,  13'd300,  -13'd176,  -13'd583,  13'd88,  -13'd241,  -13'd536,  -13'd831,  -13'd413,  13'd517,  -13'd453,  13'd10,  
13'd250,  13'd242,  -13'd310,  -13'd596,  13'd642,  -13'd599,  -13'd316,  -13'd414,  13'd421,  13'd540,  -13'd361,  13'd75,  -13'd212,  -13'd139,  -13'd396,  -13'd44,  
13'd302,  13'd55,  -13'd94,  -13'd43,  -13'd173,  -13'd109,  -13'd398,  -13'd483,  -13'd103,  13'd154,  -13'd60,  -13'd201,  -13'd389,  13'd501,  -13'd489,  -13'd95,  

13'd261,  -13'd75,  -13'd767,  -13'd605,  -13'd461,  -13'd1287,  13'd1271,  -13'd990,  13'd107,  -13'd1154,  -13'd1007,  -13'd77,  -13'd599,  13'd453,  -13'd932,  -13'd826,  
-13'd70,  13'd423,  -13'd863,  -13'd156,  -13'd176,  -13'd724,  -13'd14,  13'd27,  13'd27,  13'd534,  -13'd1040,  -13'd83,  -13'd759,  -13'd520,  -13'd141,  -13'd847,  
13'd810,  13'd508,  -13'd778,  -13'd57,  -13'd161,  13'd798,  -13'd1000,  13'd586,  -13'd123,  13'd154,  13'd165,  13'd268,  13'd77,  -13'd1518,  13'd554,  13'd477,  
13'd98,  -13'd362,  -13'd184,  13'd212,  13'd287,  13'd228,  -13'd5,  -13'd152,  13'd468,  13'd341,  13'd401,  13'd566,  13'd113,  -13'd781,  13'd351,  13'd158,  
-13'd1167,  13'd474,  13'd54,  -13'd374,  -13'd81,  13'd212,  13'd2,  -13'd429,  -13'd141,  -13'd278,  13'd365,  13'd200,  -13'd426,  13'd120,  13'd182,  13'd517,  
-13'd175,  -13'd20,  -13'd634,  13'd40,  -13'd758,  -13'd191,  13'd14,  13'd90,  -13'd420,  13'd297,  -13'd434,  -13'd31,  13'd127,  -13'd94,  -13'd442,  -13'd805,  
13'd660,  13'd300,  13'd321,  -13'd310,  13'd230,  -13'd92,  -13'd108,  13'd459,  13'd126,  -13'd190,  -13'd659,  -13'd297,  -13'd469,  -13'd60,  13'd248,  -13'd37,  
13'd235,  -13'd164,  -13'd81,  -13'd419,  -13'd666,  -13'd215,  13'd42,  13'd884,  13'd225,  13'd69,  -13'd147,  13'd115,  -13'd469,  -13'd1340,  13'd899,  -13'd255,  
13'd515,  -13'd501,  13'd40,  13'd87,  -13'd124,  13'd323,  13'd138,  13'd67,  -13'd123,  -13'd352,  -13'd446,  -13'd519,  13'd173,  13'd331,  -13'd75,  13'd95,  
-13'd872,  -13'd265,  -13'd354,  13'd276,  -13'd254,  13'd151,  13'd717,  13'd409,  13'd617,  -13'd631,  13'd819,  13'd351,  -13'd43,  13'd673,  -13'd211,  -13'd312,  
13'd616,  13'd315,  13'd740,  -13'd48,  13'd590,  -13'd74,  13'd95,  -13'd250,  -13'd228,  -13'd10,  -13'd1477,  13'd191,  -13'd168,  13'd696,  13'd152,  13'd123,  
-13'd42,  -13'd328,  13'd796,  -13'd227,  13'd455,  13'd202,  -13'd700,  13'd323,  13'd6,  13'd89,  -13'd844,  13'd266,  13'd182,  13'd358,  13'd32,  -13'd840,  
13'd112,  -13'd84,  13'd706,  13'd425,  -13'd265,  -13'd2,  13'd281,  -13'd424,  13'd33,  -13'd328,  13'd363,  -13'd152,  -13'd499,  -13'd355,  13'd183,  13'd119,  
13'd338,  13'd570,  13'd198,  -13'd769,  13'd186,  -13'd435,  -13'd122,  -13'd158,  13'd346,  13'd142,  13'd474,  -13'd609,  -13'd106,  13'd669,  -13'd472,  13'd253,  
-13'd226,  13'd2,  13'd382,  -13'd366,  13'd18,  13'd157,  13'd22,  13'd430,  13'd227,  -13'd869,  13'd391,  -13'd269,  13'd158,  13'd1082,  13'd713,  -13'd71,  
13'd60,  13'd25,  13'd449,  13'd260,  -13'd235,  -13'd82,  -13'd1173,  13'd117,  -13'd731,  13'd195,  -13'd874,  13'd37,  13'd34,  13'd358,  -13'd108,  -13'd6,  
-13'd147,  -13'd45,  13'd522,  13'd339,  -13'd47,  -13'd93,  13'd33,  -13'd91,  -13'd163,  -13'd280,  -13'd490,  13'd100,  -13'd64,  13'd256,  -13'd6,  -13'd389,  
-13'd294,  13'd1150,  13'd567,  -13'd829,  13'd607,  -13'd427,  13'd263,  -13'd247,  -13'd305,  13'd254,  -13'd17,  13'd273,  -13'd168,  -13'd76,  13'd713,  -13'd182,  
-13'd81,  13'd90,  13'd648,  -13'd8,  -13'd100,  -13'd237,  13'd516,  -13'd725,  13'd138,  -13'd670,  -13'd644,  13'd651,  13'd127,  13'd609,  -13'd834,  -13'd88,  
13'd352,  13'd681,  -13'd372,  -13'd589,  -13'd634,  -13'd16,  -13'd293,  13'd309,  -13'd372,  -13'd969,  -13'd457,  -13'd522,  13'd146,  13'd433,  -13'd968,  -13'd1166,  
-13'd669,  13'd74,  13'd416,  13'd434,  13'd1010,  13'd357,  -13'd565,  13'd36,  -13'd304,  13'd204,  13'd399,  -13'd2,  -13'd142,  -13'd37,  -13'd131,  -13'd325,  
13'd142,  13'd57,  -13'd97,  -13'd522,  13'd104,  -13'd221,  -13'd775,  -13'd208,  -13'd359,  -13'd754,  13'd297,  13'd254,  13'd257,  -13'd201,  13'd30,  13'd458,  
13'd801,  -13'd723,  -13'd180,  13'd576,  -13'd148,  -13'd101,  -13'd342,  -13'd334,  13'd735,  13'd270,  -13'd181,  13'd329,  -13'd33,  -13'd566,  -13'd161,  13'd18,  
13'd915,  -13'd207,  13'd505,  13'd243,  -13'd209,  -13'd295,  13'd192,  13'd343,  13'd300,  13'd382,  13'd49,  13'd795,  13'd180,  13'd308,  -13'd690,  13'd83,  
13'd186,  -13'd477,  -13'd718,  -13'd523,  -13'd527,  -13'd655,  -13'd147,  13'd461,  13'd934,  -13'd1053,  -13'd532,  -13'd1021,  13'd50,  13'd415,  -13'd201,  -13'd142,  

13'd122,  -13'd274,  -13'd106,  13'd12,  13'd34,  13'd523,  -13'd1158,  13'd17,  13'd225,  -13'd91,  13'd394,  -13'd516,  -13'd95,  -13'd1048,  13'd59,  -13'd244,  
-13'd56,  13'd265,  -13'd157,  13'd443,  13'd12,  -13'd278,  -13'd303,  -13'd55,  13'd929,  13'd276,  -13'd559,  -13'd831,  13'd387,  -13'd171,  -13'd192,  13'd1274,  
-13'd137,  -13'd566,  -13'd136,  -13'd707,  13'd767,  13'd68,  -13'd102,  13'd704,  13'd104,  13'd54,  -13'd926,  13'd300,  13'd305,  -13'd3,  -13'd165,  13'd287,  
-13'd722,  -13'd917,  -13'd432,  -13'd332,  13'd447,  -13'd442,  13'd138,  -13'd166,  -13'd113,  -13'd951,  -13'd391,  -13'd466,  -13'd327,  13'd1154,  -13'd548,  13'd317,  
-13'd349,  -13'd147,  13'd380,  -13'd425,  13'd436,  -13'd13,  -13'd398,  13'd54,  -13'd150,  -13'd141,  -13'd451,  13'd665,  -13'd667,  13'd336,  13'd212,  -13'd947,  
13'd159,  13'd268,  -13'd605,  -13'd322,  13'd867,  -13'd556,  -13'd381,  13'd494,  -13'd56,  -13'd530,  -13'd95,  -13'd74,  13'd48,  -13'd1147,  13'd336,  -13'd201,  
-13'd91,  13'd25,  -13'd84,  -13'd764,  13'd62,  -13'd259,  13'd340,  -13'd31,  -13'd3,  13'd462,  -13'd415,  13'd497,  -13'd380,  13'd102,  13'd374,  13'd221,  
13'd823,  -13'd406,  13'd359,  -13'd231,  13'd326,  13'd205,  13'd257,  13'd681,  -13'd71,  13'd698,  -13'd124,  13'd933,  -13'd376,  13'd709,  13'd556,  13'd447,  
13'd1207,  -13'd682,  13'd725,  13'd253,  13'd10,  13'd573,  13'd210,  13'd630,  -13'd61,  -13'd287,  13'd178,  13'd566,  -13'd105,  13'd979,  13'd295,  13'd550,  
13'd883,  13'd568,  -13'd186,  13'd16,  13'd578,  13'd452,  -13'd105,  -13'd216,  13'd52,  -13'd915,  -13'd767,  -13'd578,  13'd581,  13'd697,  -13'd241,  -13'd150,  
-13'd79,  -13'd136,  -13'd28,  13'd235,  13'd265,  13'd367,  -13'd244,  13'd317,  13'd590,  -13'd34,  13'd87,  -13'd627,  13'd196,  -13'd516,  13'd341,  13'd200,  
13'd230,  -13'd427,  -13'd448,  -13'd314,  -13'd548,  13'd353,  -13'd183,  13'd487,  13'd537,  13'd319,  13'd11,  13'd108,  13'd903,  13'd450,  -13'd21,  -13'd10,  
-13'd33,  -13'd313,  -13'd881,  13'd887,  -13'd545,  -13'd270,  -13'd52,  13'd208,  -13'd95,  13'd491,  13'd757,  13'd572,  13'd391,  -13'd713,  13'd247,  13'd679,  
-13'd68,  -13'd1125,  13'd898,  13'd368,  13'd238,  13'd168,  13'd228,  13'd812,  -13'd391,  13'd1,  13'd289,  13'd509,  13'd811,  -13'd788,  13'd172,  -13'd47,  
-13'd124,  -13'd386,  -13'd572,  -13'd165,  -13'd524,  -13'd185,  13'd632,  13'd693,  -13'd166,  13'd218,  -13'd40,  -13'd621,  13'd827,  -13'd90,  -13'd54,  13'd722,  
-13'd103,  -13'd515,  13'd676,  -13'd71,  13'd584,  -13'd35,  -13'd697,  13'd293,  13'd105,  -13'd25,  -13'd15,  -13'd10,  13'd299,  -13'd461,  -13'd45,  -13'd336,  
-13'd503,  13'd147,  13'd50,  13'd150,  13'd238,  -13'd359,  -13'd525,  13'd311,  13'd331,  -13'd255,  -13'd373,  13'd297,  13'd237,  13'd84,  -13'd9,  13'd540,  
-13'd307,  -13'd355,  -13'd516,  13'd82,  -13'd22,  -13'd403,  13'd13,  -13'd458,  -13'd489,  -13'd130,  -13'd155,  13'd113,  -13'd543,  -13'd449,  -13'd369,  13'd73,  
13'd500,  13'd678,  13'd204,  -13'd359,  -13'd1056,  13'd662,  -13'd421,  13'd26,  13'd246,  13'd251,  13'd473,  13'd199,  -13'd201,  -13'd117,  13'd211,  13'd171,  
-13'd338,  13'd134,  -13'd262,  -13'd19,  13'd757,  -13'd309,  13'd183,  13'd730,  13'd247,  -13'd525,  13'd105,  13'd495,  -13'd211,  13'd271,  13'd437,  -13'd149,  
-13'd128,  13'd163,  -13'd310,  13'd644,  13'd366,  13'd346,  -13'd294,  -13'd281,  -13'd53,  -13'd314,  -13'd126,  13'd757,  13'd174,  13'd160,  -13'd275,  -13'd308,  
13'd182,  13'd231,  -13'd725,  13'd130,  -13'd558,  -13'd445,  -13'd884,  -13'd610,  13'd164,  13'd388,  13'd239,  -13'd12,  -13'd412,  13'd236,  13'd291,  13'd253,  
-13'd35,  -13'd291,  -13'd172,  -13'd810,  13'd299,  -13'd509,  13'd448,  13'd445,  13'd322,  13'd536,  -13'd375,  13'd264,  -13'd401,  13'd606,  13'd321,  -13'd192,  
13'd170,  -13'd466,  13'd958,  -13'd293,  13'd170,  13'd168,  13'd528,  -13'd274,  13'd856,  -13'd363,  -13'd218,  13'd430,  -13'd405,  13'd157,  13'd301,  13'd83,  
13'd50,  -13'd190,  13'd402,  -13'd228,  13'd193,  -13'd309,  13'd787,  13'd625,  -13'd416,  -13'd1237,  -13'd113,  13'd494,  13'd92,  -13'd10,  -13'd242,  13'd259,  

13'd775,  13'd350,  -13'd599,  -13'd287,  -13'd354,  13'd872,  -13'd404,  13'd239,  -13'd152,  13'd45,  13'd286,  13'd253,  13'd149,  -13'd759,  13'd637,  13'd245,  
-13'd285,  13'd279,  -13'd464,  -13'd410,  -13'd345,  13'd331,  13'd323,  13'd889,  -13'd83,  13'd368,  13'd311,  13'd45,  -13'd139,  -13'd625,  13'd677,  13'd293,  
13'd98,  13'd635,  -13'd736,  13'd228,  13'd320,  13'd244,  -13'd53,  -13'd575,  -13'd338,  13'd85,  13'd53,  13'd166,  -13'd620,  13'd932,  13'd167,  13'd358,  
13'd19,  13'd131,  13'd310,  -13'd692,  -13'd159,  13'd223,  13'd216,  -13'd636,  13'd243,  13'd449,  -13'd409,  -13'd122,  -13'd33,  13'd479,  -13'd303,  -13'd406,  
-13'd250,  -13'd78,  -13'd725,  -13'd131,  13'd781,  13'd161,  -13'd350,  -13'd657,  -13'd765,  -13'd560,  -13'd110,  -13'd228,  -13'd866,  13'd531,  13'd416,  13'd554,  
13'd478,  -13'd337,  -13'd56,  13'd304,  13'd53,  -13'd440,  13'd356,  13'd323,  -13'd263,  13'd724,  13'd51,  -13'd31,  13'd336,  -13'd191,  -13'd180,  13'd569,  
13'd276,  13'd529,  -13'd149,  13'd356,  13'd415,  -13'd18,  13'd330,  -13'd666,  -13'd13,  13'd743,  -13'd651,  -13'd482,  13'd61,  13'd113,  -13'd110,  13'd768,  
-13'd147,  13'd42,  -13'd369,  -13'd297,  13'd28,  -13'd614,  -13'd606,  13'd335,  -13'd609,  13'd345,  13'd648,  13'd359,  13'd422,  -13'd393,  13'd64,  13'd541,  
13'd453,  -13'd665,  13'd124,  13'd176,  -13'd185,  -13'd210,  -13'd341,  -13'd559,  13'd98,  -13'd232,  -13'd140,  13'd85,  -13'd321,  13'd217,  -13'd583,  13'd559,  
13'd975,  13'd1061,  13'd210,  -13'd507,  -13'd82,  13'd193,  13'd292,  -13'd173,  13'd211,  -13'd297,  -13'd192,  13'd789,  13'd449,  -13'd391,  -13'd717,  -13'd649,  
-13'd479,  13'd625,  -13'd269,  -13'd209,  13'd218,  -13'd131,  -13'd200,  13'd223,  13'd85,  13'd648,  13'd449,  13'd41,  13'd80,  -13'd57,  -13'd545,  -13'd105,  
13'd566,  13'd467,  13'd421,  -13'd36,  -13'd116,  13'd400,  -13'd471,  13'd362,  13'd237,  13'd184,  -13'd57,  13'd36,  -13'd121,  -13'd298,  -13'd150,  13'd428,  
13'd705,  13'd380,  13'd312,  13'd116,  -13'd342,  13'd876,  13'd334,  13'd144,  13'd646,  -13'd105,  13'd573,  13'd341,  -13'd355,  -13'd718,  -13'd189,  13'd77,  
13'd615,  -13'd1028,  13'd153,  -13'd103,  13'd352,  13'd210,  13'd170,  -13'd277,  13'd627,  13'd456,  13'd72,  -13'd232,  -13'd201,  13'd153,  13'd713,  13'd317,  
13'd304,  13'd123,  -13'd903,  13'd540,  -13'd57,  13'd447,  -13'd20,  -13'd283,  13'd178,  13'd562,  13'd35,  -13'd77,  13'd387,  -13'd122,  -13'd65,  13'd475,  
13'd246,  -13'd102,  -13'd214,  -13'd211,  -13'd528,  13'd98,  -13'd174,  -13'd506,  13'd543,  -13'd354,  -13'd870,  13'd196,  13'd147,  13'd525,  13'd120,  -13'd462,  
13'd625,  13'd349,  13'd402,  13'd662,  13'd126,  13'd234,  13'd54,  -13'd236,  13'd407,  13'd15,  -13'd112,  -13'd79,  13'd201,  13'd859,  13'd104,  -13'd47,  
-13'd576,  13'd237,  -13'd202,  13'd393,  -13'd403,  13'd180,  13'd90,  -13'd538,  13'd860,  13'd392,  -13'd155,  -13'd175,  13'd154,  -13'd1103,  -13'd192,  13'd86,  
-13'd374,  -13'd234,  13'd85,  13'd94,  13'd66,  13'd355,  13'd216,  13'd206,  -13'd377,  13'd201,  13'd669,  -13'd343,  13'd188,  -13'd727,  13'd208,  -13'd674,  
-13'd867,  -13'd1,  -13'd320,  13'd242,  13'd178,  13'd98,  -13'd245,  -13'd280,  -13'd183,  13'd253,  13'd179,  13'd269,  13'd267,  13'd13,  -13'd59,  13'd208,  
13'd557,  -13'd142,  13'd811,  13'd464,  -13'd424,  13'd413,  -13'd16,  13'd709,  -13'd18,  13'd36,  -13'd697,  13'd404,  13'd201,  13'd751,  13'd310,  13'd21,  
13'd433,  13'd425,  13'd113,  13'd288,  13'd428,  -13'd360,  -13'd815,  13'd1071,  -13'd100,  -13'd371,  -13'd501,  -13'd29,  13'd670,  13'd563,  13'd70,  13'd7,  
-13'd882,  -13'd292,  13'd44,  13'd282,  13'd529,  13'd223,  13'd175,  13'd22,  -13'd1114,  -13'd1744,  13'd177,  13'd147,  13'd416,  -13'd694,  13'd191,  -13'd377,  
-13'd699,  13'd245,  -13'd731,  -13'd177,  -13'd438,  -13'd5,  -13'd182,  13'd175,  13'd385,  -13'd802,  13'd56,  13'd408,  -13'd189,  -13'd21,  13'd513,  -13'd521,  
-13'd340,  13'd359,  13'd238,  13'd395,  -13'd184,  -13'd106,  13'd325,  -13'd98,  13'd23,  -13'd521,  13'd355,  13'd541,  13'd233,  -13'd189,  -13'd125,  13'd38,  

13'd452,  13'd398,  13'd169,  13'd298,  -13'd1068,  13'd337,  13'd1227,  -13'd28,  13'd185,  -13'd520,  -13'd779,  13'd577,  -13'd970,  13'd92,  -13'd450,  13'd89,  
13'd119,  13'd80,  -13'd435,  -13'd704,  -13'd434,  13'd326,  -13'd467,  -13'd531,  13'd378,  13'd131,  13'd1005,  -13'd160,  -13'd630,  13'd601,  -13'd521,  -13'd313,  
13'd210,  13'd133,  -13'd1087,  -13'd280,  13'd435,  13'd155,  -13'd473,  -13'd481,  -13'd349,  13'd381,  13'd189,  -13'd401,  -13'd423,  13'd557,  -13'd431,  13'd539,  
-13'd374,  13'd358,  13'd6,  13'd384,  13'd492,  -13'd183,  -13'd305,  -13'd217,  13'd240,  13'd248,  -13'd62,  -13'd114,  13'd93,  13'd51,  -13'd158,  -13'd217,  
13'd345,  13'd1230,  13'd340,  -13'd347,  13'd199,  13'd434,  -13'd182,  13'd533,  -13'd337,  13'd129,  13'd193,  13'd321,  13'd597,  13'd189,  13'd403,  13'd536,  
13'd236,  -13'd160,  13'd227,  -13'd90,  13'd64,  13'd425,  -13'd252,  -13'd23,  -13'd203,  13'd317,  -13'd492,  13'd371,  -13'd60,  13'd1378,  -13'd272,  13'd267,  
13'd385,  -13'd155,  13'd281,  13'd309,  -13'd563,  13'd82,  -13'd154,  13'd492,  13'd130,  13'd184,  -13'd419,  -13'd670,  13'd793,  13'd688,  13'd831,  -13'd38,  
-13'd945,  -13'd536,  13'd108,  -13'd713,  -13'd298,  -13'd456,  -13'd260,  -13'd85,  13'd428,  13'd37,  13'd520,  -13'd2,  -13'd451,  -13'd233,  13'd118,  -13'd298,  
-13'd1007,  -13'd379,  -13'd111,  -13'd429,  -13'd211,  13'd782,  -13'd607,  13'd371,  -13'd8,  -13'd63,  -13'd279,  13'd503,  -13'd94,  -13'd140,  13'd290,  -13'd349,  
-13'd277,  13'd572,  -13'd482,  -13'd109,  13'd357,  13'd240,  13'd280,  13'd195,  13'd435,  13'd464,  -13'd416,  -13'd439,  -13'd313,  13'd146,  -13'd125,  13'd94,  
13'd446,  13'd210,  -13'd134,  13'd893,  13'd204,  13'd1366,  -13'd1141,  13'd684,  -13'd747,  13'd491,  -13'd435,  13'd510,  13'd454,  13'd298,  13'd448,  13'd489,  
-13'd397,  13'd1019,  13'd290,  13'd456,  13'd541,  -13'd318,  -13'd937,  13'd642,  13'd44,  -13'd507,  13'd1046,  13'd694,  -13'd402,  13'd186,  13'd28,  13'd820,  
-13'd469,  -13'd315,  13'd244,  13'd442,  13'd70,  13'd351,  -13'd356,  13'd779,  13'd728,  -13'd1229,  13'd263,  -13'd162,  13'd191,  -13'd8,  13'd133,  -13'd33,  
-13'd166,  13'd18,  -13'd652,  13'd80,  -13'd752,  13'd9,  -13'd96,  -13'd30,  13'd322,  13'd40,  13'd16,  13'd177,  13'd120,  -13'd89,  -13'd581,  13'd427,  
13'd171,  13'd40,  -13'd624,  -13'd39,  13'd85,  13'd53,  -13'd779,  13'd166,  -13'd403,  13'd94,  -13'd53,  -13'd115,  13'd228,  13'd55,  13'd44,  13'd391,  
13'd727,  13'd585,  -13'd145,  -13'd114,  13'd763,  -13'd108,  -13'd725,  13'd526,  -13'd276,  -13'd113,  -13'd597,  13'd518,  13'd400,  13'd564,  -13'd37,  13'd476,  
13'd149,  13'd840,  13'd769,  -13'd272,  13'd583,  13'd662,  13'd336,  -13'd320,  -13'd359,  13'd313,  -13'd45,  -13'd160,  -13'd748,  13'd228,  13'd93,  13'd367,  
13'd71,  13'd188,  13'd93,  -13'd45,  13'd170,  13'd108,  13'd423,  -13'd304,  13'd1079,  -13'd32,  -13'd324,  -13'd171,  -13'd515,  -13'd461,  -13'd300,  13'd375,  
-13'd703,  13'd592,  -13'd373,  -13'd311,  13'd443,  -13'd258,  13'd155,  13'd205,  -13'd346,  13'd176,  13'd48,  -13'd80,  -13'd603,  13'd363,  -13'd209,  -13'd268,  
-13'd327,  -13'd597,  13'd443,  -13'd148,  13'd201,  -13'd177,  13'd0,  -13'd465,  -13'd832,  -13'd13,  13'd390,  13'd91,  -13'd428,  13'd24,  -13'd248,  -13'd2,  
13'd809,  -13'd152,  13'd84,  13'd117,  -13'd30,  -13'd367,  13'd306,  13'd305,  13'd601,  -13'd421,  -13'd517,  13'd42,  13'd203,  13'd58,  13'd56,  -13'd72,  
-13'd546,  -13'd308,  13'd0,  13'd47,  13'd32,  -13'd238,  -13'd626,  13'd179,  -13'd136,  13'd414,  -13'd5,  -13'd413,  -13'd176,  -13'd21,  -13'd108,  -13'd10,  
-13'd298,  -13'd272,  13'd312,  13'd116,  -13'd364,  -13'd308,  -13'd664,  13'd203,  -13'd106,  13'd205,  -13'd432,  -13'd91,  -13'd178,  -13'd280,  13'd346,  13'd210,  
-13'd620,  13'd256,  -13'd134,  13'd723,  -13'd118,  13'd396,  -13'd143,  -13'd151,  -13'd182,  -13'd432,  13'd14,  13'd493,  -13'd34,  13'd792,  13'd102,  -13'd239,  
-13'd407,  -13'd483,  -13'd131,  13'd466,  -13'd389,  -13'd367,  -13'd3,  -13'd154,  13'd81,  -13'd834,  -13'd416,  13'd295,  13'd175,  -13'd213,  13'd115,  13'd736,  

-13'd171,  13'd36,  13'd17,  -13'd55,  13'd297,  -13'd174,  -13'd774,  13'd581,  -13'd47,  13'd188,  -13'd969,  -13'd440,  13'd496,  -13'd12,  -13'd799,  -13'd59,  
-13'd666,  13'd266,  13'd730,  13'd337,  13'd710,  -13'd32,  -13'd871,  -13'd450,  -13'd193,  13'd516,  -13'd562,  13'd268,  13'd298,  13'd677,  13'd609,  13'd748,  
13'd71,  -13'd530,  13'd256,  -13'd435,  13'd67,  -13'd437,  -13'd76,  13'd115,  13'd38,  -13'd303,  13'd70,  13'd646,  -13'd246,  13'd782,  13'd548,  13'd634,  
13'd58,  -13'd227,  13'd546,  13'd286,  -13'd19,  13'd207,  13'd408,  13'd390,  -13'd116,  -13'd139,  13'd77,  13'd502,  -13'd446,  13'd1044,  13'd652,  -13'd122,  
13'd615,  -13'd464,  13'd31,  -13'd223,  -13'd422,  -13'd336,  13'd616,  -13'd345,  13'd503,  -13'd19,  -13'd120,  13'd268,  -13'd422,  13'd228,  13'd300,  -13'd337,  
-13'd252,  -13'd451,  13'd224,  -13'd56,  13'd266,  13'd245,  -13'd768,  13'd517,  -13'd769,  13'd153,  -13'd528,  -13'd139,  -13'd222,  13'd425,  13'd118,  -13'd594,  
13'd429,  13'd432,  13'd380,  13'd749,  -13'd86,  13'd438,  13'd189,  -13'd146,  13'd236,  13'd8,  13'd442,  13'd857,  -13'd354,  13'd2,  13'd361,  -13'd654,  
-13'd197,  13'd496,  13'd666,  13'd353,  13'd170,  13'd230,  13'd319,  13'd713,  13'd536,  13'd47,  13'd98,  -13'd217,  13'd28,  13'd1057,  13'd422,  -13'd715,  
-13'd430,  13'd302,  13'd236,  13'd173,  -13'd271,  13'd158,  13'd236,  13'd311,  -13'd177,  -13'd973,  13'd517,  13'd397,  -13'd736,  13'd80,  13'd256,  -13'd54,  
13'd365,  13'd461,  13'd22,  -13'd484,  13'd368,  13'd142,  13'd280,  -13'd339,  13'd416,  -13'd662,  -13'd54,  -13'd333,  13'd62,  -13'd827,  13'd293,  13'd443,  
13'd642,  13'd5,  -13'd188,  -13'd189,  13'd143,  -13'd485,  -13'd131,  -13'd176,  13'd720,  13'd129,  13'd1273,  -13'd340,  -13'd370,  13'd496,  13'd115,  -13'd49,  
13'd64,  13'd540,  13'd178,  -13'd303,  -13'd526,  13'd384,  13'd96,  13'd733,  -13'd332,  13'd148,  13'd299,  -13'd54,  13'd127,  13'd58,  13'd110,  13'd636,  
13'd200,  13'd429,  13'd324,  13'd299,  13'd179,  -13'd178,  13'd133,  13'd447,  -13'd303,  13'd96,  13'd10,  13'd392,  13'd183,  13'd707,  -13'd100,  -13'd251,  
-13'd543,  13'd142,  13'd483,  -13'd25,  -13'd10,  13'd40,  13'd634,  13'd38,  -13'd213,  -13'd226,  13'd685,  13'd185,  -13'd342,  -13'd347,  -13'd239,  -13'd928,  
13'd335,  13'd8,  -13'd250,  13'd298,  13'd308,  13'd190,  13'd234,  13'd102,  -13'd36,  -13'd1417,  -13'd431,  -13'd653,  -13'd275,  13'd50,  13'd238,  -13'd682,  
-13'd75,  13'd427,  -13'd171,  -13'd199,  13'd1153,  -13'd505,  -13'd719,  13'd54,  13'd619,  -13'd389,  13'd201,  -13'd146,  13'd167,  13'd49,  -13'd854,  13'd77,  
-13'd224,  -13'd631,  -13'd143,  13'd287,  -13'd27,  -13'd36,  13'd537,  -13'd157,  -13'd212,  -13'd195,  13'd284,  13'd215,  -13'd23,  13'd251,  -13'd437,  13'd351,  
13'd579,  -13'd171,  -13'd52,  13'd136,  -13'd232,  13'd899,  -13'd115,  -13'd593,  13'd221,  13'd31,  13'd191,  -13'd609,  13'd346,  13'd405,  13'd201,  -13'd122,  
-13'd27,  -13'd486,  -13'd24,  13'd174,  13'd462,  -13'd818,  -13'd514,  -13'd2,  13'd1059,  13'd132,  13'd271,  -13'd260,  -13'd477,  13'd61,  13'd6,  13'd517,  
13'd576,  -13'd108,  13'd162,  -13'd399,  -13'd313,  -13'd336,  -13'd378,  -13'd42,  -13'd19,  13'd255,  -13'd471,  13'd167,  13'd235,  -13'd288,  -13'd265,  -13'd54,  
-13'd581,  -13'd350,  -13'd866,  -13'd146,  -13'd408,  13'd38,  -13'd50,  13'd158,  13'd408,  -13'd382,  13'd1017,  -13'd16,  -13'd211,  13'd156,  13'd70,  13'd183,  
-13'd88,  13'd330,  -13'd676,  13'd9,  -13'd250,  13'd380,  13'd432,  -13'd1021,  13'd778,  -13'd597,  13'd281,  13'd835,  -13'd621,  13'd211,  13'd17,  13'd233,  
-13'd129,  13'd501,  13'd196,  -13'd753,  -13'd33,  -13'd37,  13'd532,  -13'd354,  13'd426,  13'd614,  13'd227,  -13'd30,  13'd115,  13'd853,  13'd107,  13'd736,  
13'd282,  -13'd25,  13'd670,  13'd552,  -13'd143,  -13'd470,  -13'd221,  -13'd209,  -13'd480,  13'd274,  -13'd516,  -13'd353,  -13'd780,  13'd246,  13'd377,  -13'd254,  
13'd831,  13'd740,  13'd804,  -13'd212,  13'd624,  13'd703,  -13'd456,  13'd172,  -13'd106,  13'd1152,  -13'd488,  13'd431,  -13'd182,  13'd495,  13'd218,  13'd178,  

13'd615,  -13'd48,  13'd229,  13'd252,  13'd559,  -13'd163,  13'd369,  13'd193,  13'd317,  13'd72,  -13'd260,  -13'd100,  13'd338,  -13'd483,  13'd191,  13'd251,  
-13'd374,  -13'd164,  13'd255,  -13'd239,  -13'd498,  -13'd187,  13'd1199,  13'd392,  13'd131,  -13'd471,  13'd511,  -13'd475,  -13'd142,  13'd284,  -13'd762,  -13'd258,  
-13'd42,  13'd547,  -13'd154,  13'd244,  13'd231,  -13'd8,  -13'd114,  13'd400,  13'd63,  -13'd258,  13'd50,  -13'd359,  -13'd491,  -13'd714,  -13'd104,  -13'd277,  
13'd604,  13'd660,  13'd293,  13'd438,  -13'd284,  -13'd483,  -13'd279,  -13'd170,  -13'd9,  13'd162,  13'd199,  13'd399,  13'd1018,  -13'd1042,  -13'd4,  -13'd518,  
13'd723,  13'd812,  -13'd555,  13'd482,  -13'd221,  -13'd32,  -13'd57,  -13'd150,  -13'd359,  13'd697,  -13'd444,  13'd263,  13'd408,  13'd341,  -13'd472,  13'd221,  
-13'd333,  -13'd333,  13'd319,  -13'd624,  -13'd208,  -13'd575,  -13'd121,  -13'd65,  13'd452,  -13'd146,  13'd798,  -13'd114,  13'd311,  -13'd123,  13'd227,  -13'd499,  
-13'd277,  -13'd736,  13'd175,  13'd569,  13'd119,  -13'd390,  13'd342,  13'd448,  13'd399,  -13'd605,  13'd352,  13'd684,  13'd203,  13'd682,  13'd363,  -13'd780,  
13'd189,  -13'd558,  13'd234,  13'd442,  -13'd488,  -13'd495,  -13'd603,  13'd82,  13'd558,  -13'd588,  13'd823,  -13'd598,  13'd234,  -13'd88,  13'd156,  13'd142,  
-13'd899,  13'd286,  -13'd839,  13'd249,  13'd335,  -13'd581,  -13'd557,  13'd634,  13'd247,  13'd1150,  13'd302,  13'd111,  13'd752,  -13'd796,  13'd409,  13'd537,  
-13'd289,  -13'd450,  -13'd107,  13'd422,  13'd485,  13'd372,  -13'd709,  -13'd106,  -13'd794,  13'd1635,  13'd477,  -13'd48,  -13'd97,  -13'd468,  13'd199,  13'd447,  
-13'd224,  13'd165,  -13'd174,  13'd284,  -13'd1061,  13'd103,  13'd198,  -13'd336,  -13'd118,  -13'd362,  -13'd749,  -13'd773,  -13'd349,  13'd750,  13'd9,  13'd189,  
13'd150,  -13'd152,  -13'd448,  13'd93,  -13'd376,  13'd301,  -13'd6,  13'd403,  -13'd193,  13'd34,  -13'd618,  -13'd755,  13'd154,  -13'd74,  13'd109,  13'd519,  
-13'd929,  13'd554,  -13'd754,  13'd178,  13'd272,  -13'd225,  13'd349,  13'd418,  13'd897,  13'd505,  13'd20,  -13'd343,  -13'd393,  -13'd321,  13'd534,  13'd620,  
-13'd1004,  13'd174,  -13'd1092,  -13'd201,  13'd553,  -13'd25,  -13'd180,  13'd182,  -13'd108,  13'd419,  13'd578,  13'd456,  -13'd415,  -13'd224,  -13'd34,  13'd807,  
-13'd270,  -13'd368,  13'd852,  -13'd26,  13'd491,  13'd581,  13'd665,  13'd537,  13'd747,  13'd384,  13'd111,  13'd987,  -13'd102,  -13'd183,  13'd86,  -13'd227,  
13'd290,  -13'd170,  -13'd105,  13'd103,  -13'd138,  13'd273,  13'd81,  13'd409,  13'd306,  -13'd107,  -13'd504,  -13'd333,  -13'd398,  -13'd98,  -13'd433,  13'd307,  
-13'd496,  -13'd24,  -13'd58,  -13'd136,  -13'd439,  13'd375,  13'd192,  13'd766,  -13'd765,  -13'd62,  13'd216,  13'd288,  -13'd69,  13'd57,  13'd444,  -13'd342,  
13'd16,  -13'd819,  -13'd293,  -13'd94,  13'd478,  13'd132,  13'd49,  13'd354,  -13'd546,  -13'd402,  13'd632,  13'd728,  13'd577,  -13'd64,  13'd8,  13'd5,  
13'd266,  13'd938,  -13'd223,  -13'd63,  13'd89,  13'd951,  -13'd461,  -13'd521,  13'd719,  -13'd580,  13'd195,  -13'd251,  13'd526,  13'd314,  13'd35,  -13'd439,  
-13'd68,  -13'd94,  13'd942,  13'd14,  -13'd156,  13'd119,  13'd299,  13'd1,  -13'd249,  -13'd449,  13'd752,  -13'd410,  -13'd304,  13'd523,  13'd183,  13'd50,  
13'd290,  -13'd367,  -13'd553,  -13'd61,  -13'd254,  13'd717,  -13'd249,  -13'd264,  -13'd135,  13'd219,  -13'd9,  13'd88,  -13'd810,  13'd311,  13'd510,  -13'd17,  
-13'd274,  13'd26,  -13'd380,  13'd435,  -13'd263,  13'd885,  13'd259,  -13'd170,  13'd73,  13'd528,  13'd90,  13'd249,  13'd65,  -13'd1026,  -13'd145,  -13'd110,  
13'd539,  13'd170,  -13'd793,  -13'd289,  -13'd73,  13'd282,  13'd643,  -13'd667,  -13'd185,  -13'd98,  13'd886,  -13'd80,  -13'd100,  -13'd771,  13'd229,  13'd100,  
-13'd327,  13'd402,  13'd206,  -13'd487,  13'd241,  -13'd397,  13'd859,  -13'd170,  13'd486,  -13'd249,  -13'd98,  -13'd484,  -13'd405,  13'd746,  13'd119,  -13'd79,  
-13'd289,  -13'd150,  -13'd427,  -13'd621,  -13'd461,  13'd90,  -13'd265,  -13'd232,  13'd796,  13'd59,  -13'd479,  -13'd621,  13'd125,  13'd39,  -13'd1073,  13'd41,  

-13'd140,  -13'd287,  13'd66,  13'd213,  -13'd288,  13'd276,  13'd127,  13'd290,  -13'd340,  13'd229,  -13'd804,  -13'd880,  13'd167,  13'd204,  -13'd51,  13'd43,  
-13'd852,  13'd18,  13'd307,  -13'd88,  -13'd15,  -13'd362,  -13'd152,  -13'd224,  -13'd525,  -13'd536,  -13'd525,  -13'd367,  -13'd855,  13'd609,  13'd383,  13'd134,  
-13'd68,  -13'd213,  13'd474,  -13'd22,  -13'd363,  13'd548,  -13'd846,  13'd387,  13'd699,  -13'd541,  13'd616,  13'd320,  13'd41,  13'd1018,  13'd177,  -13'd264,  
-13'd372,  13'd897,  13'd780,  -13'd362,  -13'd195,  -13'd148,  13'd332,  13'd522,  13'd262,  -13'd142,  13'd122,  -13'd314,  -13'd49,  -13'd1123,  13'd453,  13'd583,  
-13'd532,  -13'd526,  -13'd43,  13'd387,  -13'd220,  -13'd931,  -13'd186,  -13'd417,  13'd375,  13'd105,  -13'd22,  -13'd68,  -13'd431,  13'd100,  13'd467,  -13'd807,  
-13'd27,  13'd207,  -13'd848,  13'd9,  13'd340,  13'd254,  -13'd896,  -13'd745,  -13'd250,  13'd108,  -13'd297,  -13'd110,  -13'd136,  -13'd1019,  -13'd449,  -13'd639,  
13'd716,  -13'd343,  13'd180,  13'd849,  -13'd328,  -13'd198,  13'd415,  -13'd75,  -13'd913,  13'd409,  13'd336,  -13'd26,  -13'd145,  -13'd396,  -13'd562,  -13'd381,  
13'd175,  -13'd90,  13'd369,  -13'd671,  -13'd778,  -13'd53,  13'd497,  13'd97,  -13'd214,  13'd861,  13'd132,  13'd485,  13'd309,  -13'd83,  -13'd522,  13'd59,  
-13'd154,  -13'd249,  13'd345,  -13'd200,  -13'd609,  -13'd124,  -13'd63,  13'd391,  -13'd581,  13'd21,  -13'd380,  13'd74,  -13'd65,  -13'd185,  13'd382,  -13'd90,  
-13'd1111,  13'd513,  13'd866,  -13'd161,  -13'd495,  -13'd908,  -13'd163,  -13'd252,  -13'd105,  13'd595,  13'd311,  13'd132,  -13'd416,  13'd84,  13'd221,  13'd250,  
-13'd199,  13'd58,  -13'd829,  13'd308,  -13'd81,  -13'd361,  -13'd539,  13'd53,  13'd964,  13'd118,  13'd1044,  13'd26,  -13'd209,  -13'd867,  13'd129,  13'd493,  
13'd641,  -13'd603,  -13'd925,  13'd343,  -13'd233,  13'd435,  -13'd222,  13'd305,  13'd365,  13'd903,  13'd256,  13'd694,  13'd552,  -13'd1248,  -13'd186,  13'd429,  
13'd902,  -13'd268,  13'd177,  13'd591,  13'd819,  -13'd443,  13'd411,  13'd719,  13'd1018,  13'd566,  13'd300,  13'd206,  13'd894,  -13'd364,  13'd75,  13'd94,  
-13'd56,  -13'd634,  -13'd220,  13'd441,  -13'd67,  13'd310,  -13'd47,  -13'd272,  13'd360,  13'd666,  -13'd331,  13'd34,  -13'd465,  13'd1253,  -13'd6,  -13'd256,  
13'd1645,  13'd655,  13'd1030,  13'd215,  -13'd1356,  13'd448,  -13'd232,  13'd195,  13'd393,  -13'd159,  -13'd386,  13'd66,  13'd875,  -13'd587,  13'd281,  -13'd224,  
13'd351,  -13'd667,  13'd149,  -13'd3,  13'd1,  -13'd529,  13'd934,  -13'd226,  13'd1575,  13'd672,  13'd880,  -13'd180,  13'd193,  13'd398,  13'd245,  13'd367,  
-13'd318,  -13'd219,  -13'd247,  13'd20,  -13'd85,  13'd336,  -13'd8,  13'd330,  13'd249,  -13'd114,  13'd1324,  13'd416,  13'd590,  13'd546,  13'd528,  -13'd61,  
-13'd621,  13'd559,  -13'd95,  13'd849,  13'd122,  13'd638,  13'd209,  -13'd328,  -13'd709,  -13'd713,  13'd583,  13'd113,  13'd171,  -13'd58,  13'd651,  13'd229,  
-13'd359,  13'd101,  -13'd643,  -13'd51,  13'd307,  -13'd571,  13'd196,  13'd16,  -13'd346,  13'd440,  -13'd529,  -13'd1080,  13'd647,  13'd12,  13'd146,  -13'd591,  
13'd860,  -13'd320,  13'd946,  -13'd610,  13'd715,  -13'd749,  -13'd566,  13'd447,  13'd23,  13'd606,  13'd702,  13'd28,  13'd310,  13'd253,  -13'd628,  -13'd138,  
13'd1,  -13'd219,  -13'd339,  -13'd8,  -13'd199,  13'd264,  13'd521,  13'd293,  -13'd285,  -13'd308,  13'd106,  -13'd972,  13'd706,  13'd222,  13'd29,  13'd240,  
-13'd937,  13'd96,  -13'd760,  13'd30,  -13'd494,  -13'd510,  13'd262,  -13'd552,  -13'd153,  -13'd454,  13'd251,  -13'd691,  13'd504,  13'd257,  13'd126,  13'd351,  
-13'd702,  -13'd285,  -13'd305,  -13'd314,  -13'd406,  -13'd35,  -13'd574,  13'd100,  -13'd912,  -13'd379,  13'd119,  -13'd708,  -13'd890,  13'd250,  -13'd472,  13'd750,  
-13'd666,  13'd168,  -13'd1167,  13'd240,  -13'd67,  -13'd64,  -13'd170,  13'd98,  13'd23,  -13'd460,  13'd263,  13'd300,  -13'd430,  -13'd837,  13'd156,  -13'd140,  
-13'd1541,  13'd619,  -13'd621,  -13'd124,  -13'd348,  -13'd967,  -13'd307,  -13'd237,  -13'd821,  13'd79,  13'd343,  -13'd157,  -13'd678,  13'd357,  -13'd437,  -13'd320,  

13'd94,  -13'd56,  13'd361,  -13'd51,  13'd338,  -13'd271,  -13'd377,  13'd678,  13'd211,  13'd426,  13'd113,  13'd913,  13'd96,  13'd911,  13'd135,  13'd412,  
13'd164,  -13'd268,  13'd227,  13'd165,  13'd60,  13'd403,  13'd572,  13'd246,  13'd534,  -13'd120,  13'd713,  13'd682,  13'd441,  13'd541,  -13'd19,  13'd12,  
13'd587,  13'd197,  -13'd393,  -13'd585,  -13'd929,  -13'd147,  -13'd234,  13'd96,  13'd339,  13'd16,  -13'd95,  13'd51,  13'd579,  13'd388,  -13'd666,  -13'd612,  
13'd485,  13'd403,  -13'd862,  13'd309,  -13'd307,  13'd47,  13'd382,  13'd254,  -13'd541,  13'd19,  13'd594,  -13'd104,  13'd132,  13'd160,  -13'd322,  13'd627,  
13'd807,  13'd1208,  -13'd741,  -13'd394,  13'd641,  13'd334,  13'd256,  -13'd136,  -13'd206,  13'd311,  13'd394,  13'd64,  13'd1138,  -13'd46,  13'd64,  13'd167,  
-13'd420,  13'd775,  13'd101,  13'd53,  13'd552,  13'd861,  -13'd255,  -13'd285,  13'd289,  13'd20,  -13'd335,  13'd901,  13'd13,  13'd644,  13'd313,  13'd285,  
13'd138,  13'd49,  13'd233,  13'd824,  13'd198,  -13'd378,  13'd85,  -13'd254,  -13'd342,  13'd23,  13'd736,  13'd262,  13'd112,  -13'd61,  13'd189,  -13'd355,  
-13'd962,  -13'd534,  13'd209,  13'd120,  -13'd355,  13'd367,  13'd393,  -13'd4,  13'd720,  -13'd749,  -13'd26,  -13'd473,  13'd362,  -13'd501,  13'd116,  13'd138,  
-13'd284,  13'd238,  -13'd133,  13'd85,  13'd49,  -13'd619,  -13'd605,  -13'd684,  13'd439,  13'd376,  13'd81,  13'd425,  -13'd113,  -13'd197,  -13'd202,  13'd515,  
13'd27,  -13'd944,  -13'd169,  13'd574,  13'd1005,  13'd637,  -13'd70,  13'd108,  -13'd95,  -13'd18,  -13'd475,  -13'd6,  13'd489,  -13'd1112,  -13'd479,  13'd816,  
-13'd266,  13'd160,  13'd73,  13'd8,  13'd732,  -13'd100,  13'd211,  -13'd488,  13'd38,  13'd294,  13'd557,  13'd213,  13'd271,  -13'd415,  -13'd108,  13'd687,  
-13'd113,  13'd255,  13'd443,  13'd456,  13'd280,  13'd468,  13'd456,  -13'd61,  -13'd509,  -13'd426,  13'd287,  -13'd126,  -13'd25,  -13'd107,  13'd359,  -13'd337,  
13'd67,  -13'd713,  13'd163,  -13'd363,  -13'd45,  13'd83,  13'd429,  -13'd573,  13'd97,  -13'd324,  -13'd149,  13'd49,  -13'd546,  -13'd262,  -13'd316,  -13'd298,  
-13'd581,  -13'd596,  -13'd965,  13'd199,  -13'd56,  -13'd224,  13'd41,  -13'd521,  13'd399,  -13'd188,  -13'd138,  13'd36,  13'd77,  -13'd58,  13'd480,  -13'd30,  
-13'd369,  -13'd395,  -13'd406,  -13'd41,  13'd270,  13'd128,  -13'd37,  13'd38,  -13'd450,  13'd737,  13'd823,  13'd93,  13'd285,  13'd636,  13'd648,  13'd653,  
13'd37,  13'd329,  13'd21,  -13'd741,  -13'd730,  -13'd152,  13'd441,  -13'd513,  -13'd363,  13'd150,  -13'd445,  13'd119,  -13'd174,  -13'd290,  -13'd261,  13'd545,  
13'd995,  13'd84,  13'd39,  13'd309,  13'd619,  -13'd599,  13'd105,  -13'd451,  -13'd816,  13'd46,  -13'd780,  13'd174,  13'd296,  13'd464,  13'd375,  -13'd61,  
13'd163,  13'd798,  13'd409,  -13'd100,  13'd511,  -13'd27,  13'd452,  -13'd388,  13'd556,  -13'd190,  13'd741,  -13'd710,  -13'd301,  -13'd680,  13'd195,  -13'd16,  
13'd53,  -13'd125,  -13'd617,  13'd728,  -13'd146,  13'd92,  13'd105,  -13'd803,  -13'd204,  13'd739,  -13'd266,  -13'd272,  -13'd93,  -13'd636,  13'd339,  13'd61,  
-13'd832,  -13'd140,  13'd638,  13'd488,  13'd162,  -13'd459,  -13'd36,  13'd238,  -13'd367,  13'd365,  -13'd172,  13'd780,  -13'd317,  13'd487,  -13'd641,  13'd63,  
13'd360,  -13'd75,  -13'd624,  -13'd80,  -13'd371,  -13'd292,  -13'd884,  -13'd530,  -13'd622,  13'd643,  -13'd134,  13'd26,  13'd41,  13'd1290,  -13'd523,  -13'd199,  
13'd15,  13'd418,  -13'd421,  13'd128,  -13'd217,  -13'd195,  -13'd996,  -13'd13,  13'd233,  -13'd321,  -13'd545,  -13'd375,  13'd29,  13'd184,  13'd172,  -13'd287,  
13'd477,  -13'd76,  -13'd1006,  -13'd264,  -13'd277,  13'd457,  -13'd25,  13'd528,  -13'd277,  -13'd902,  13'd521,  -13'd251,  -13'd303,  -13'd352,  13'd372,  13'd317,  
13'd535,  13'd338,  -13'd255,  13'd317,  -13'd308,  13'd60,  -13'd290,  13'd387,  13'd32,  -13'd797,  13'd71,  13'd214,  13'd216,  -13'd27,  -13'd113,  13'd127,  
-13'd640,  -13'd315,  -13'd793,  -13'd234,  -13'd217,  -13'd271,  13'd124,  13'd134,  -13'd783,  -13'd1671,  -13'd334,  -13'd853,  -13'd651,  -13'd79,  -13'd76,  -13'd447,  

13'd444,  13'd404,  13'd899,  13'd629,  13'd424,  13'd157,  13'd551,  13'd275,  13'd631,  13'd454,  13'd289,  -13'd347,  13'd323,  13'd959,  13'd545,  -13'd775,  
-13'd727,  -13'd740,  13'd532,  13'd539,  13'd488,  -13'd3,  -13'd310,  -13'd335,  -13'd254,  13'd597,  13'd125,  13'd162,  -13'd63,  -13'd80,  -13'd64,  13'd87,  
-13'd307,  -13'd32,  -13'd53,  13'd149,  -13'd351,  13'd313,  13'd138,  13'd296,  13'd24,  13'd94,  13'd547,  13'd802,  13'd103,  -13'd1260,  -13'd241,  -13'd832,  
13'd399,  -13'd49,  -13'd72,  -13'd144,  13'd817,  -13'd627,  -13'd654,  13'd77,  -13'd443,  13'd570,  -13'd33,  -13'd460,  13'd622,  -13'd1352,  -13'd842,  13'd589,  
13'd767,  -13'd872,  -13'd769,  -13'd24,  -13'd496,  13'd59,  -13'd547,  13'd752,  -13'd175,  13'd181,  -13'd256,  -13'd824,  -13'd126,  -13'd466,  -13'd182,  -13'd238,  
-13'd355,  13'd565,  -13'd583,  13'd568,  13'd457,  13'd203,  -13'd506,  13'd627,  13'd282,  13'd299,  13'd644,  13'd135,  -13'd153,  -13'd50,  13'd872,  -13'd179,  
-13'd187,  -13'd231,  13'd265,  13'd369,  13'd303,  13'd279,  13'd89,  13'd325,  13'd253,  13'd426,  13'd201,  13'd396,  -13'd343,  -13'd575,  -13'd264,  -13'd434,  
-13'd1329,  13'd484,  -13'd775,  -13'd291,  13'd625,  -13'd763,  13'd525,  13'd600,  -13'd63,  13'd21,  13'd269,  13'd159,  13'd118,  -13'd155,  13'd194,  -13'd85,  
13'd305,  13'd22,  -13'd10,  13'd363,  13'd185,  -13'd42,  -13'd762,  -13'd92,  -13'd496,  13'd150,  13'd4,  -13'd6,  13'd302,  -13'd6,  13'd209,  -13'd40,  
13'd953,  -13'd224,  -13'd917,  -13'd17,  -13'd371,  13'd6,  -13'd430,  13'd18,  13'd45,  13'd726,  13'd327,  13'd211,  13'd546,  -13'd981,  13'd262,  13'd547,  
13'd323,  13'd85,  -13'd177,  13'd191,  13'd852,  -13'd348,  -13'd223,  13'd84,  -13'd369,  -13'd844,  13'd411,  13'd180,  13'd102,  -13'd18,  -13'd122,  -13'd217,  
-13'd9,  13'd60,  -13'd115,  -13'd484,  -13'd508,  -13'd272,  -13'd459,  -13'd738,  -13'd137,  -13'd15,  13'd805,  -13'd103,  13'd37,  -13'd770,  13'd537,  13'd198,  
13'd68,  -13'd365,  13'd277,  13'd240,  -13'd492,  -13'd245,  -13'd232,  13'd310,  -13'd76,  -13'd518,  13'd1368,  -13'd515,  -13'd253,  13'd655,  13'd717,  13'd244,  
-13'd63,  13'd421,  13'd106,  13'd546,  13'd114,  13'd26,  13'd135,  -13'd2,  13'd576,  -13'd649,  13'd132,  13'd212,  13'd622,  -13'd226,  -13'd142,  13'd382,  
-13'd1227,  -13'd450,  13'd356,  13'd895,  13'd252,  13'd336,  13'd13,  -13'd215,  13'd209,  13'd260,  13'd438,  13'd130,  13'd763,  13'd115,  13'd708,  -13'd166,  
13'd386,  13'd268,  13'd156,  -13'd283,  13'd209,  -13'd478,  13'd120,  13'd231,  -13'd541,  -13'd57,  13'd613,  13'd29,  13'd381,  -13'd259,  13'd29,  -13'd133,  
-13'd396,  13'd71,  -13'd852,  -13'd628,  -13'd104,  -13'd970,  -13'd83,  -13'd292,  -13'd165,  -13'd152,  13'd266,  13'd123,  13'd135,  13'd103,  -13'd908,  13'd361,  
13'd578,  13'd749,  13'd7,  -13'd822,  13'd133,  -13'd679,  13'd167,  -13'd50,  13'd195,  13'd417,  -13'd22,  -13'd288,  -13'd207,  13'd639,  -13'd62,  -13'd45,  
13'd691,  13'd907,  13'd823,  -13'd578,  -13'd5,  -13'd133,  13'd143,  13'd601,  13'd752,  13'd277,  13'd320,  13'd605,  -13'd620,  -13'd52,  13'd736,  -13'd410,  
13'd138,  13'd355,  -13'd57,  13'd526,  13'd688,  13'd228,  -13'd86,  13'd117,  13'd258,  -13'd60,  13'd670,  -13'd727,  13'd69,  13'd367,  -13'd268,  13'd621,  
-13'd21,  13'd85,  -13'd211,  -13'd881,  13'd24,  -13'd273,  13'd433,  -13'd818,  13'd163,  -13'd1043,  -13'd687,  13'd293,  -13'd1030,  -13'd793,  13'd103,  13'd341,  
-13'd280,  -13'd171,  -13'd900,  -13'd67,  -13'd26,  -13'd103,  13'd636,  -13'd394,  13'd798,  -13'd385,  -13'd506,  13'd263,  -13'd351,  13'd151,  -13'd205,  13'd31,  
13'd509,  -13'd316,  13'd610,  -13'd243,  13'd378,  -13'd105,  13'd677,  -13'd634,  13'd1548,  13'd183,  -13'd96,  -13'd52,  -13'd446,  13'd526,  -13'd231,  -13'd561,  
-13'd296,  13'd173,  13'd316,  -13'd354,  -13'd10,  -13'd322,  -13'd406,  13'd431,  13'd13,  13'd16,  -13'd472,  -13'd393,  -13'd32,  13'd668,  13'd74,  -13'd277,  
-13'd421,  13'd118,  13'd213,  13'd233,  -13'd476,  13'd117,  -13'd420,  -13'd41,  13'd198,  13'd947,  13'd132,  -13'd166,  -13'd615,  -13'd211,  -13'd733,  -13'd175,  

13'd198,  13'd918,  13'd251,  -13'd208,  -13'd362,  13'd52,  13'd1161,  -13'd283,  13'd53,  -13'd58,  -13'd68,  13'd1064,  -13'd860,  13'd797,  -13'd814,  13'd162,  
13'd10,  13'd380,  -13'd398,  -13'd224,  -13'd828,  -13'd312,  13'd994,  13'd112,  13'd549,  -13'd165,  -13'd98,  13'd85,  -13'd615,  13'd2,  13'd176,  13'd137,  
13'd861,  13'd305,  -13'd14,  -13'd579,  13'd418,  -13'd498,  -13'd194,  13'd307,  13'd531,  -13'd6,  13'd39,  13'd27,  13'd194,  13'd46,  13'd23,  -13'd260,  
-13'd37,  -13'd114,  13'd44,  13'd168,  -13'd54,  13'd679,  13'd261,  13'd22,  13'd266,  13'd268,  -13'd200,  -13'd343,  13'd488,  -13'd369,  -13'd128,  -13'd2,  
-13'd1077,  13'd752,  13'd395,  -13'd141,  -13'd538,  13'd539,  -13'd259,  13'd27,  13'd219,  -13'd154,  13'd725,  13'd36,  13'd531,  13'd776,  13'd618,  13'd685,  
-13'd580,  -13'd718,  13'd131,  -13'd552,  -13'd401,  -13'd209,  13'd581,  13'd160,  13'd510,  -13'd243,  -13'd71,  -13'd196,  -13'd703,  13'd187,  13'd259,  13'd153,  
13'd446,  -13'd169,  13'd215,  -13'd774,  13'd203,  13'd64,  -13'd582,  -13'd309,  13'd458,  13'd222,  -13'd318,  -13'd226,  -13'd187,  13'd591,  13'd397,  13'd32,  
-13'd574,  -13'd438,  -13'd19,  -13'd431,  13'd228,  -13'd267,  13'd120,  13'd526,  -13'd312,  13'd352,  13'd538,  13'd290,  -13'd853,  -13'd277,  13'd87,  -13'd400,  
-13'd140,  -13'd29,  -13'd34,  -13'd268,  13'd449,  13'd94,  -13'd150,  -13'd318,  -13'd438,  13'd1136,  -13'd190,  -13'd28,  13'd44,  -13'd504,  13'd67,  -13'd119,  
-13'd642,  -13'd574,  -13'd163,  -13'd163,  -13'd541,  -13'd725,  13'd406,  13'd143,  13'd59,  13'd251,  -13'd302,  -13'd213,  -13'd320,  -13'd279,  -13'd857,  13'd415,  
-13'd329,  13'd490,  -13'd146,  -13'd45,  13'd157,  13'd682,  -13'd361,  13'd148,  -13'd759,  13'd821,  -13'd522,  -13'd138,  13'd70,  -13'd34,  13'd198,  13'd108,  
13'd947,  13'd376,  13'd142,  13'd78,  -13'd47,  13'd214,  -13'd2,  13'd490,  -13'd69,  -13'd163,  13'd267,  -13'd425,  -13'd949,  13'd835,  13'd128,  -13'd721,  
-13'd213,  13'd472,  -13'd431,  -13'd38,  13'd773,  13'd286,  13'd170,  13'd300,  13'd752,  -13'd361,  -13'd197,  13'd682,  -13'd398,  -13'd454,  -13'd339,  -13'd577,  
13'd144,  13'd136,  -13'd558,  -13'd1217,  13'd449,  13'd389,  13'd230,  -13'd558,  13'd829,  13'd542,  -13'd203,  -13'd536,  13'd61,  -13'd54,  -13'd129,  -13'd147,  
-13'd664,  -13'd411,  -13'd392,  13'd595,  -13'd835,  13'd527,  -13'd511,  -13'd157,  13'd401,  13'd543,  13'd194,  -13'd52,  -13'd870,  -13'd78,  -13'd75,  13'd771,  
13'd105,  -13'd97,  13'd748,  13'd382,  -13'd78,  13'd154,  -13'd68,  -13'd137,  -13'd366,  -13'd156,  -13'd885,  13'd555,  -13'd288,  13'd244,  -13'd12,  13'd362,  
13'd593,  13'd178,  -13'd383,  13'd655,  -13'd134,  13'd209,  -13'd399,  13'd108,  13'd942,  -13'd353,  -13'd603,  13'd351,  13'd442,  13'd305,  13'd787,  13'd288,  
-13'd332,  -13'd317,  -13'd38,  13'd63,  -13'd91,  13'd177,  13'd663,  13'd781,  -13'd577,  -13'd593,  13'd8,  -13'd154,  -13'd947,  13'd388,  13'd462,  -13'd126,  
-13'd38,  13'd305,  -13'd272,  13'd79,  13'd422,  13'd311,  -13'd149,  -13'd726,  -13'd270,  -13'd107,  -13'd427,  13'd547,  -13'd29,  13'd998,  13'd42,  -13'd374,  
-13'd358,  13'd269,  13'd644,  13'd253,  -13'd204,  13'd321,  13'd583,  -13'd476,  13'd642,  13'd96,  -13'd207,  -13'd22,  -13'd514,  13'd485,  -13'd206,  -13'd77,  
-13'd813,  -13'd563,  -13'd304,  13'd493,  13'd370,  13'd1009,  -13'd363,  13'd974,  13'd298,  13'd147,  -13'd394,  -13'd437,  13'd510,  -13'd576,  13'd32,  13'd327,  
13'd28,  13'd587,  13'd86,  13'd373,  13'd1134,  -13'd7,  -13'd507,  13'd1033,  -13'd333,  -13'd547,  13'd896,  -13'd451,  -13'd13,  -13'd411,  13'd679,  -13'd18,  
-13'd345,  -13'd350,  -13'd418,  13'd610,  13'd63,  13'd618,  -13'd197,  13'd669,  13'd222,  13'd560,  13'd534,  13'd97,  13'd498,  -13'd104,  13'd37,  13'd252,  
13'd43,  13'd712,  -13'd547,  13'd830,  -13'd208,  13'd795,  13'd2,  13'd352,  13'd129,  13'd571,  -13'd531,  13'd1048,  13'd677,  -13'd60,  13'd64,  -13'd260,  
13'd977,  13'd221,  13'd327,  13'd758,  13'd299,  13'd145,  13'd257,  13'd862,  13'd1391,  13'd216,  13'd361,  13'd699,  -13'd25,  13'd486,  -13'd155,  -13'd160,  

-13'd158,  -13'd84,  13'd173,  13'd72,  -13'd83,  13'd232,  13'd706,  13'd492,  -13'd629,  -13'd383,  -13'd122,  -13'd61,  -13'd187,  -13'd576,  13'd83,  -13'd160,  
13'd99,  -13'd638,  13'd66,  -13'd553,  13'd172,  -13'd108,  -13'd517,  -13'd865,  -13'd815,  -13'd421,  -13'd252,  -13'd561,  13'd75,  13'd121,  -13'd803,  -13'd615,  
-13'd32,  13'd118,  13'd232,  13'd375,  -13'd597,  -13'd209,  -13'd363,  -13'd117,  -13'd39,  13'd89,  -13'd65,  -13'd960,  13'd41,  13'd337,  -13'd545,  13'd421,  
-13'd638,  -13'd304,  -13'd622,  13'd137,  13'd244,  -13'd772,  -13'd86,  -13'd294,  13'd149,  -13'd377,  -13'd174,  13'd87,  -13'd93,  13'd29,  -13'd132,  -13'd61,  
-13'd43,  13'd120,  -13'd468,  -13'd404,  13'd8,  -13'd146,  -13'd146,  13'd66,  13'd133,  13'd487,  -13'd343,  13'd65,  13'd123,  -13'd331,  -13'd516,  -13'd516,  
-13'd325,  -13'd295,  -13'd187,  -13'd324,  -13'd768,  13'd524,  -13'd498,  13'd450,  13'd457,  -13'd21,  -13'd365,  -13'd547,  13'd496,  -13'd236,  13'd399,  -13'd581,  
-13'd32,  13'd53,  13'd21,  13'd446,  13'd337,  13'd520,  -13'd543,  -13'd907,  -13'd137,  13'd547,  13'd483,  -13'd227,  13'd301,  13'd300,  13'd302,  -13'd607,  
13'd560,  13'd351,  -13'd332,  -13'd685,  13'd190,  13'd301,  -13'd95,  13'd124,  -13'd218,  -13'd40,  -13'd522,  13'd203,  13'd209,  13'd294,  -13'd397,  -13'd531,  
-13'd270,  -13'd95,  -13'd514,  13'd1,  13'd65,  -13'd452,  -13'd597,  -13'd539,  -13'd198,  13'd142,  -13'd493,  -13'd170,  -13'd544,  -13'd163,  13'd185,  -13'd253,  
13'd545,  13'd226,  13'd687,  -13'd419,  -13'd369,  13'd323,  -13'd229,  -13'd221,  -13'd404,  13'd276,  -13'd235,  -13'd661,  -13'd609,  13'd301,  -13'd507,  13'd171,  
-13'd377,  -13'd535,  -13'd588,  13'd119,  -13'd317,  13'd215,  -13'd308,  -13'd815,  13'd388,  -13'd396,  -13'd823,  -13'd133,  -13'd168,  -13'd141,  -13'd140,  -13'd420,  
13'd176,  -13'd387,  -13'd31,  -13'd195,  -13'd653,  -13'd149,  13'd182,  -13'd375,  -13'd381,  13'd338,  -13'd295,  -13'd487,  -13'd498,  -13'd308,  13'd242,  -13'd421,  
13'd214,  -13'd110,  -13'd709,  13'd227,  -13'd277,  -13'd792,  -13'd19,  13'd255,  -13'd153,  -13'd365,  13'd122,  -13'd850,  -13'd319,  -13'd194,  13'd413,  -13'd28,  
13'd176,  -13'd545,  -13'd731,  13'd611,  -13'd348,  -13'd70,  -13'd76,  -13'd318,  -13'd789,  13'd9,  -13'd453,  -13'd616,  -13'd265,  -13'd123,  13'd444,  -13'd120,  
13'd252,  13'd167,  -13'd480,  13'd168,  -13'd11,  -13'd181,  -13'd385,  -13'd66,  -13'd460,  13'd414,  -13'd225,  -13'd190,  13'd106,  13'd688,  -13'd275,  13'd510,  
-13'd6,  13'd209,  -13'd443,  -13'd346,  -13'd129,  -13'd171,  13'd126,  -13'd196,  13'd233,  -13'd498,  13'd372,  -13'd261,  -13'd420,  13'd3,  -13'd226,  -13'd96,  
13'd433,  -13'd454,  13'd245,  -13'd16,  -13'd625,  -13'd552,  -13'd132,  13'd77,  -13'd24,  -13'd792,  -13'd268,  13'd203,  -13'd14,  -13'd241,  -13'd926,  -13'd288,  
13'd464,  -13'd254,  -13'd564,  -13'd410,  13'd289,  -13'd358,  -13'd290,  -13'd270,  13'd131,  -13'd823,  -13'd430,  -13'd141,  13'd260,  -13'd860,  13'd339,  13'd167,  
13'd20,  -13'd295,  13'd168,  -13'd191,  -13'd52,  13'd487,  13'd288,  -13'd466,  -13'd391,  13'd180,  -13'd249,  13'd33,  13'd80,  -13'd242,  -13'd693,  -13'd388,  
13'd52,  -13'd202,  -13'd411,  -13'd837,  13'd234,  13'd245,  -13'd835,  -13'd874,  -13'd43,  13'd356,  -13'd83,  13'd346,  -13'd680,  -13'd23,  13'd11,  13'd98,  
-13'd280,  -13'd456,  -13'd898,  -13'd230,  -13'd721,  -13'd776,  -13'd150,  -13'd746,  -13'd581,  -13'd425,  -13'd86,  -13'd169,  -13'd293,  13'd401,  -13'd319,  -13'd104,  
-13'd482,  13'd74,  -13'd143,  -13'd818,  -13'd584,  -13'd582,  13'd106,  -13'd618,  13'd288,  -13'd295,  -13'd473,  13'd126,  -13'd437,  -13'd267,  -13'd834,  13'd15,  
13'd508,  -13'd171,  -13'd117,  13'd187,  -13'd37,  -13'd84,  -13'd358,  13'd82,  13'd344,  13'd19,  -13'd223,  -13'd715,  -13'd56,  -13'd529,  13'd30,  -13'd36,  
13'd652,  13'd252,  13'd405,  -13'd770,  -13'd168,  13'd73,  -13'd535,  -13'd278,  -13'd609,  13'd328,  -13'd771,  13'd105,  -13'd748,  13'd315,  -13'd638,  -13'd246,  
13'd682,  13'd524,  -13'd84,  -13'd478,  -13'd180,  -13'd505,  13'd164,  -13'd22,  13'd235,  -13'd22,  13'd611,  -13'd546,  -13'd171,  13'd45,  -13'd15,  -13'd523,  

13'd295,  -13'd684,  13'd368,  -13'd299,  -13'd526,  -13'd102,  -13'd418,  -13'd328,  -13'd62,  13'd883,  -13'd739,  -13'd758,  -13'd771,  -13'd322,  -13'd977,  -13'd201,  
-13'd520,  -13'd1143,  -13'd309,  -13'd25,  -13'd137,  13'd615,  13'd65,  -13'd3,  -13'd1111,  -13'd1,  -13'd624,  -13'd923,  -13'd592,  -13'd1114,  -13'd540,  13'd113,  
-13'd219,  13'd300,  -13'd25,  13'd334,  -13'd692,  13'd246,  -13'd1182,  -13'd264,  -13'd204,  -13'd456,  -13'd1036,  13'd281,  -13'd241,  13'd135,  -13'd884,  -13'd394,  
-13'd138,  13'd391,  -13'd20,  13'd61,  13'd114,  13'd946,  -13'd246,  -13'd622,  13'd332,  -13'd213,  -13'd619,  -13'd591,  -13'd498,  -13'd749,  -13'd163,  13'd218,  
13'd887,  13'd647,  13'd351,  13'd672,  -13'd547,  13'd382,  -13'd254,  13'd377,  13'd431,  -13'd327,  -13'd128,  -13'd654,  -13'd309,  -13'd277,  13'd112,  13'd233,  
-13'd738,  -13'd480,  -13'd1052,  13'd105,  -13'd285,  -13'd516,  -13'd1093,  -13'd731,  -13'd209,  13'd354,  13'd917,  13'd744,  13'd104,  -13'd136,  -13'd135,  -13'd603,  
-13'd275,  -13'd356,  13'd97,  13'd423,  13'd88,  13'd373,  -13'd307,  -13'd507,  13'd437,  13'd372,  13'd962,  -13'd532,  13'd368,  -13'd94,  -13'd57,  -13'd0,  
13'd506,  13'd215,  13'd198,  13'd522,  13'd75,  13'd264,  -13'd55,  13'd885,  13'd116,  13'd434,  -13'd5,  -13'd81,  13'd817,  13'd690,  13'd168,  -13'd107,  
13'd1017,  13'd11,  -13'd93,  -13'd134,  13'd269,  13'd710,  -13'd331,  13'd141,  13'd803,  -13'd104,  13'd1270,  -13'd299,  13'd371,  13'd492,  -13'd127,  -13'd2,  
13'd228,  13'd268,  13'd298,  -13'd136,  13'd821,  -13'd682,  -13'd706,  -13'd55,  -13'd268,  13'd1085,  -13'd787,  13'd512,  -13'd306,  13'd927,  13'd0,  13'd241,  
-13'd681,  13'd110,  -13'd879,  13'd79,  -13'd247,  13'd443,  13'd723,  13'd252,  13'd1198,  -13'd189,  13'd843,  -13'd597,  -13'd41,  13'd350,  13'd712,  13'd609,  
-13'd336,  13'd42,  -13'd273,  13'd170,  -13'd55,  -13'd300,  13'd204,  -13'd614,  13'd720,  -13'd50,  13'd486,  -13'd474,  -13'd920,  13'd962,  13'd829,  13'd546,  
-13'd211,  -13'd377,  -13'd350,  -13'd519,  13'd56,  -13'd954,  -13'd428,  13'd275,  -13'd916,  -13'd210,  -13'd322,  -13'd925,  -13'd110,  13'd230,  13'd742,  13'd573,  
13'd217,  13'd324,  -13'd530,  -13'd215,  -13'd385,  -13'd589,  -13'd1052,  -13'd162,  -13'd518,  -13'd186,  13'd20,  -13'd421,  -13'd964,  13'd668,  13'd179,  13'd138,  
13'd523,  -13'd167,  13'd803,  -13'd352,  -13'd394,  -13'd577,  13'd74,  -13'd813,  13'd294,  13'd931,  -13'd818,  13'd824,  -13'd638,  13'd198,  13'd194,  13'd337,  
-13'd134,  -13'd934,  13'd618,  -13'd75,  -13'd305,  -13'd378,  13'd101,  -13'd233,  -13'd645,  13'd78,  13'd893,  -13'd688,  -13'd709,  -13'd705,  -13'd680,  -13'd58,  
13'd243,  -13'd360,  -13'd435,  13'd313,  -13'd507,  -13'd705,  -13'd284,  13'd105,  -13'd842,  -13'd773,  13'd179,  -13'd838,  -13'd40,  -13'd156,  -13'd516,  13'd127,  
13'd94,  13'd777,  -13'd230,  -13'd54,  -13'd570,  -13'd329,  13'd399,  13'd277,  13'd1011,  13'd501,  -13'd540,  -13'd476,  -13'd845,  -13'd310,  -13'd385,  -13'd612,  
13'd228,  13'd477,  13'd102,  -13'd421,  -13'd881,  13'd139,  13'd48,  13'd292,  13'd293,  13'd27,  13'd61,  13'd352,  -13'd447,  13'd254,  -13'd144,  -13'd491,  
13'd778,  -13'd235,  13'd238,  -13'd121,  -13'd667,  13'd603,  13'd221,  13'd511,  13'd402,  -13'd90,  13'd452,  13'd80,  13'd626,  13'd425,  13'd644,  13'd232,  
-13'd781,  13'd856,  -13'd992,  -13'd764,  13'd564,  -13'd608,  -13'd916,  -13'd782,  -13'd306,  -13'd743,  -13'd460,  13'd327,  -13'd162,  13'd365,  -13'd320,  -13'd152,  
-13'd170,  13'd343,  13'd170,  -13'd1212,  -13'd158,  -13'd554,  -13'd428,  -13'd747,  -13'd710,  -13'd331,  13'd174,  -13'd110,  -13'd584,  13'd159,  -13'd14,  -13'd648,  
13'd584,  -13'd398,  13'd680,  -13'd57,  -13'd578,  -13'd365,  -13'd483,  -13'd107,  13'd687,  -13'd114,  -13'd1136,  -13'd14,  -13'd949,  13'd62,  13'd278,  -13'd675,  
13'd942,  -13'd887,  13'd520,  13'd13,  13'd531,  13'd157,  -13'd301,  -13'd510,  13'd39,  13'd711,  13'd292,  -13'd12,  13'd158,  13'd114,  13'd149,  -13'd18,  
13'd584,  -13'd341,  -13'd742,  -13'd139,  13'd136,  13'd561,  -13'd30,  13'd516,  13'd343,  -13'd2,  13'd311,  13'd314,  -13'd34,  -13'd350,  13'd1061,  13'd538,  

-13'd133,  -13'd587,  -13'd263,  13'd922,  13'd182,  13'd666,  13'd308,  13'd588,  13'd467,  13'd344,  13'd816,  -13'd14,  13'd426,  -13'd288,  13'd294,  -13'd9,  
-13'd807,  -13'd404,  13'd690,  13'd855,  13'd81,  13'd416,  -13'd328,  13'd544,  13'd208,  13'd961,  13'd698,  -13'd615,  13'd573,  -13'd241,  13'd979,  -13'd373,  
-13'd414,  -13'd908,  -13'd205,  -13'd2,  -13'd635,  13'd125,  -13'd436,  13'd485,  -13'd63,  13'd121,  -13'd108,  13'd170,  13'd695,  -13'd1493,  -13'd217,  -13'd153,  
13'd384,  13'd182,  -13'd88,  13'd338,  13'd303,  13'd276,  -13'd378,  -13'd274,  -13'd317,  13'd53,  -13'd455,  13'd378,  13'd755,  -13'd1510,  -13'd303,  -13'd102,  
-13'd35,  13'd157,  13'd90,  13'd131,  -13'd277,  13'd204,  -13'd254,  -13'd123,  -13'd471,  -13'd466,  -13'd581,  -13'd165,  13'd939,  -13'd153,  -13'd55,  13'd291,  
-13'd327,  -13'd426,  -13'd330,  13'd275,  -13'd194,  -13'd280,  -13'd1033,  13'd129,  -13'd208,  -13'd262,  13'd494,  13'd6,  13'd60,  13'd692,  13'd180,  -13'd96,  
-13'd148,  13'd170,  -13'd186,  13'd246,  13'd12,  13'd98,  -13'd85,  -13'd106,  13'd449,  -13'd673,  13'd181,  13'd250,  13'd340,  13'd377,  -13'd114,  -13'd267,  
-13'd970,  13'd443,  -13'd195,  13'd176,  -13'd466,  13'd345,  -13'd781,  -13'd284,  13'd1409,  13'd91,  13'd356,  13'd85,  13'd74,  -13'd614,  -13'd152,  13'd357,  
-13'd63,  -13'd266,  -13'd689,  -13'd143,  -13'd473,  -13'd418,  -13'd831,  13'd422,  13'd425,  13'd808,  -13'd279,  13'd289,  13'd873,  -13'd1163,  -13'd306,  13'd519,  
13'd258,  13'd101,  -13'd500,  -13'd100,  13'd783,  13'd130,  13'd252,  13'd257,  13'd444,  13'd300,  13'd547,  -13'd299,  13'd101,  -13'd194,  -13'd744,  13'd264,  
-13'd237,  -13'd20,  13'd606,  13'd174,  -13'd342,  13'd301,  -13'd82,  13'd409,  13'd1,  -13'd89,  -13'd159,  -13'd647,  13'd206,  13'd209,  -13'd682,  13'd194,  
13'd178,  13'd6,  13'd762,  -13'd259,  -13'd160,  -13'd394,  13'd573,  13'd241,  -13'd341,  -13'd685,  13'd470,  -13'd420,  -13'd297,  -13'd320,  13'd393,  13'd236,  
13'd325,  13'd156,  13'd282,  -13'd373,  -13'd515,  -13'd187,  13'd277,  -13'd183,  -13'd369,  13'd100,  -13'd77,  -13'd626,  -13'd18,  13'd36,  -13'd116,  13'd870,  
-13'd529,  13'd624,  -13'd92,  13'd130,  13'd88,  13'd645,  -13'd76,  13'd413,  13'd523,  13'd36,  -13'd177,  -13'd239,  13'd241,  -13'd67,  13'd248,  13'd500,  
-13'd1574,  -13'd196,  -13'd511,  -13'd166,  -13'd56,  -13'd899,  13'd181,  13'd50,  13'd119,  -13'd113,  13'd829,  13'd394,  -13'd532,  -13'd223,  13'd772,  13'd233,  
13'd138,  -13'd69,  13'd14,  -13'd149,  -13'd577,  -13'd312,  13'd571,  -13'd852,  13'd453,  -13'd23,  13'd215,  -13'd196,  -13'd113,  13'd93,  -13'd735,  -13'd770,  
-13'd315,  -13'd280,  -13'd361,  -13'd487,  -13'd234,  13'd132,  -13'd282,  13'd419,  -13'd679,  13'd1021,  13'd712,  13'd324,  -13'd254,  13'd1,  -13'd2,  13'd93,  
-13'd52,  13'd188,  -13'd362,  13'd339,  13'd140,  13'd4,  -13'd601,  13'd464,  13'd438,  -13'd500,  -13'd400,  -13'd212,  13'd133,  13'd553,  -13'd8,  -13'd725,  
13'd150,  -13'd82,  13'd615,  -13'd104,  13'd215,  13'd184,  -13'd1,  -13'd179,  -13'd509,  -13'd410,  13'd465,  13'd25,  -13'd549,  -13'd113,  -13'd531,  -13'd383,  
13'd326,  13'd601,  13'd483,  -13'd363,  -13'd40,  -13'd140,  13'd377,  13'd544,  13'd94,  -13'd17,  13'd240,  -13'd20,  -13'd218,  13'd609,  -13'd113,  -13'd673,  
13'd294,  -13'd160,  -13'd102,  13'd649,  -13'd566,  -13'd627,  13'd921,  13'd30,  13'd962,  13'd270,  13'd265,  13'd95,  -13'd324,  -13'd1003,  13'd29,  13'd526,  
-13'd248,  13'd14,  -13'd726,  13'd562,  -13'd211,  13'd165,  13'd444,  -13'd145,  13'd211,  -13'd332,  13'd14,  -13'd149,  -13'd320,  13'd231,  -13'd604,  13'd461,  
13'd352,  -13'd163,  13'd579,  -13'd584,  -13'd85,  -13'd392,  -13'd107,  13'd224,  13'd1113,  -13'd104,  13'd351,  13'd90,  -13'd162,  13'd109,  -13'd740,  -13'd436,  
13'd234,  13'd680,  13'd114,  13'd285,  -13'd330,  -13'd174,  -13'd47,  -13'd72,  13'd889,  -13'd70,  13'd312,  -13'd543,  13'd259,  13'd203,  -13'd47,  -13'd102,  
13'd143,  13'd317,  -13'd101,  -13'd922,  -13'd596,  -13'd524,  -13'd130,  -13'd61,  -13'd31,  -13'd475,  -13'd467,  -13'd501,  -13'd213,  13'd414,  -13'd204,  -13'd240,  

-13'd692,  13'd238,  13'd601,  13'd811,  13'd53,  13'd263,  -13'd1192,  13'd1185,  -13'd247,  13'd1106,  -13'd998,  13'd120,  13'd484,  -13'd410,  -13'd120,  -13'd41,  
-13'd28,  13'd476,  13'd1745,  13'd278,  13'd657,  -13'd67,  -13'd91,  13'd540,  13'd560,  -13'd25,  -13'd421,  -13'd193,  -13'd177,  13'd967,  -13'd276,  -13'd772,  
13'd347,  13'd145,  13'd1483,  13'd347,  -13'd701,  13'd201,  13'd522,  -13'd306,  13'd116,  -13'd492,  -13'd102,  -13'd144,  -13'd305,  13'd1021,  13'd400,  -13'd655,  
13'd104,  -13'd4,  13'd142,  13'd615,  -13'd158,  -13'd515,  13'd254,  13'd239,  -13'd415,  -13'd9,  13'd721,  13'd441,  13'd561,  -13'd349,  -13'd488,  -13'd517,  
13'd542,  13'd1073,  -13'd430,  -13'd52,  -13'd337,  13'd782,  13'd259,  -13'd188,  13'd491,  13'd247,  13'd539,  -13'd381,  13'd598,  13'd437,  -13'd186,  13'd335,  
-13'd186,  13'd841,  13'd894,  13'd28,  13'd667,  13'd813,  -13'd775,  13'd127,  -13'd281,  13'd88,  -13'd535,  -13'd135,  13'd519,  13'd345,  13'd151,  13'd416,  
13'd592,  13'd153,  13'd697,  13'd597,  -13'd139,  13'd483,  -13'd378,  -13'd81,  13'd815,  -13'd86,  -13'd312,  13'd276,  -13'd173,  13'd407,  13'd54,  -13'd68,  
13'd398,  13'd354,  13'd1183,  13'd688,  -13'd267,  13'd2,  -13'd601,  13'd126,  -13'd197,  -13'd10,  13'd498,  -13'd313,  -13'd765,  13'd743,  13'd282,  -13'd234,  
13'd19,  13'd573,  13'd1005,  -13'd652,  -13'd348,  13'd51,  13'd67,  -13'd172,  -13'd135,  -13'd362,  -13'd413,  13'd101,  13'd186,  13'd379,  -13'd376,  -13'd270,  
13'd253,  13'd124,  -13'd531,  13'd562,  13'd8,  -13'd810,  -13'd134,  -13'd191,  13'd311,  -13'd305,  13'd824,  -13'd343,  -13'd169,  13'd113,  -13'd473,  13'd15,  
-13'd603,  13'd165,  -13'd538,  13'd497,  13'd390,  13'd176,  -13'd249,  13'd601,  13'd426,  13'd280,  13'd761,  13'd323,  13'd440,  13'd15,  13'd246,  13'd290,  
-13'd99,  -13'd400,  -13'd3,  13'd344,  13'd662,  -13'd66,  13'd659,  -13'd150,  13'd619,  13'd73,  -13'd496,  -13'd417,  13'd173,  -13'd59,  13'd498,  13'd538,  
-13'd399,  13'd322,  13'd975,  -13'd364,  -13'd136,  13'd87,  -13'd358,  13'd442,  -13'd161,  -13'd467,  -13'd97,  13'd162,  -13'd57,  13'd481,  -13'd278,  -13'd318,  
-13'd800,  -13'd388,  -13'd860,  13'd503,  -13'd99,  -13'd228,  -13'd201,  13'd439,  -13'd281,  13'd314,  13'd483,  -13'd6,  -13'd635,  -13'd400,  13'd446,  13'd27,  
-13'd901,  13'd81,  13'd724,  13'd306,  -13'd29,  -13'd622,  -13'd53,  13'd115,  -13'd485,  13'd199,  13'd557,  -13'd988,  -13'd294,  -13'd769,  13'd676,  -13'd284,  
-13'd709,  13'd204,  -13'd235,  -13'd168,  -13'd167,  -13'd70,  -13'd240,  -13'd692,  13'd228,  13'd219,  13'd845,  -13'd167,  -13'd18,  -13'd564,  -13'd371,  -13'd75,  
13'd97,  -13'd121,  13'd41,  -13'd0,  13'd353,  13'd179,  -13'd324,  -13'd38,  -13'd126,  13'd1029,  -13'd553,  -13'd247,  -13'd231,  13'd410,  -13'd479,  -13'd85,  
-13'd951,  13'd62,  13'd175,  -13'd146,  13'd209,  -13'd451,  -13'd545,  13'd161,  -13'd490,  13'd216,  -13'd902,  -13'd141,  13'd360,  13'd704,  13'd546,  -13'd443,  
-13'd553,  13'd114,  13'd7,  -13'd184,  -13'd819,  -13'd117,  13'd558,  -13'd495,  -13'd191,  -13'd304,  13'd263,  13'd399,  -13'd692,  -13'd706,  -13'd157,  -13'd17,  
13'd376,  13'd401,  13'd1046,  -13'd798,  13'd87,  13'd600,  -13'd211,  13'd294,  -13'd200,  13'd213,  13'd480,  13'd962,  -13'd84,  13'd152,  -13'd534,  -13'd98,  
-13'd456,  -13'd240,  -13'd349,  -13'd614,  -13'd217,  13'd146,  13'd107,  -13'd57,  -13'd129,  13'd381,  -13'd449,  -13'd606,  -13'd494,  -13'd261,  -13'd167,  13'd283,  
-13'd149,  -13'd482,  13'd148,  13'd51,  -13'd172,  -13'd144,  -13'd336,  -13'd23,  -13'd446,  13'd79,  13'd151,  -13'd594,  -13'd79,  13'd1380,  13'd684,  13'd362,  
-13'd334,  13'd143,  13'd737,  -13'd69,  -13'd531,  13'd476,  -13'd336,  -13'd451,  -13'd462,  -13'd481,  -13'd624,  -13'd65,  -13'd271,  -13'd50,  13'd239,  -13'd252,  
13'd562,  13'd545,  13'd182,  -13'd407,  13'd432,  -13'd571,  -13'd37,  -13'd310,  -13'd401,  -13'd703,  13'd1011,  -13'd316,  -13'd171,  -13'd54,  -13'd85,  13'd348,  
13'd429,  -13'd185,  -13'd274,  13'd205,  13'd589,  13'd404,  13'd135,  -13'd239,  13'd54,  -13'd943,  -13'd175,  13'd615,  -13'd134,  13'd544,  13'd252,  13'd45,  

13'd255,  13'd819,  13'd439,  -13'd42,  -13'd247,  13'd828,  -13'd1287,  13'd435,  13'd647,  13'd229,  13'd217,  -13'd1005,  13'd654,  -13'd68,  -13'd41,  13'd633,  
-13'd246,  13'd1012,  13'd842,  13'd206,  13'd274,  -13'd115,  -13'd5,  13'd543,  13'd497,  -13'd556,  13'd655,  13'd190,  -13'd221,  13'd19,  13'd914,  -13'd190,  
-13'd24,  13'd140,  13'd142,  -13'd193,  -13'd310,  13'd87,  -13'd97,  -13'd345,  13'd242,  -13'd654,  13'd7,  -13'd2,  -13'd125,  13'd169,  13'd730,  13'd580,  
-13'd279,  -13'd202,  -13'd90,  13'd150,  -13'd844,  13'd1135,  13'd266,  13'd474,  -13'd117,  -13'd419,  13'd995,  13'd88,  13'd233,  13'd594,  13'd553,  -13'd303,  
13'd680,  13'd143,  13'd3,  -13'd104,  -13'd845,  13'd534,  13'd59,  -13'd319,  -13'd62,  -13'd740,  -13'd78,  -13'd320,  13'd168,  13'd375,  -13'd680,  13'd43,  
-13'd858,  13'd478,  13'd208,  -13'd1093,  13'd943,  -13'd236,  13'd914,  -13'd57,  -13'd49,  13'd507,  -13'd1,  -13'd466,  13'd80,  -13'd210,  -13'd447,  -13'd141,  
-13'd547,  -13'd400,  -13'd182,  -13'd1080,  13'd334,  13'd835,  -13'd432,  13'd62,  -13'd245,  -13'd322,  -13'd972,  -13'd529,  13'd161,  13'd335,  -13'd288,  -13'd433,  
13'd224,  -13'd215,  13'd468,  -13'd172,  -13'd867,  -13'd806,  -13'd708,  -13'd655,  -13'd747,  13'd133,  -13'd13,  -13'd27,  -13'd623,  -13'd93,  13'd154,  -13'd402,  
-13'd144,  -13'd63,  -13'd64,  -13'd477,  -13'd928,  13'd344,  -13'd130,  -13'd368,  -13'd31,  -13'd223,  13'd49,  -13'd568,  -13'd816,  13'd210,  -13'd30,  -13'd859,  
-13'd920,  -13'd626,  13'd1053,  13'd60,  -13'd599,  -13'd444,  -13'd36,  13'd349,  -13'd630,  13'd186,  13'd77,  -13'd410,  -13'd662,  13'd162,  13'd158,  13'd325,  
-13'd305,  -13'd454,  -13'd431,  -13'd241,  -13'd396,  -13'd355,  13'd243,  13'd289,  13'd781,  -13'd149,  -13'd878,  -13'd520,  -13'd577,  -13'd76,  13'd9,  -13'd204,  
-13'd308,  -13'd647,  13'd45,  13'd641,  -13'd205,  -13'd66,  13'd337,  -13'd547,  -13'd118,  13'd42,  -13'd925,  13'd490,  -13'd43,  -13'd85,  13'd300,  -13'd774,  
13'd54,  -13'd63,  13'd869,  13'd119,  13'd334,  -13'd449,  -13'd494,  -13'd144,  13'd1067,  -13'd84,  13'd71,  13'd1028,  -13'd119,  13'd1005,  -13'd928,  13'd182,  
-13'd776,  -13'd393,  -13'd1191,  13'd410,  -13'd56,  13'd169,  13'd217,  -13'd403,  -13'd435,  -13'd663,  13'd699,  13'd329,  13'd133,  13'd515,  -13'd734,  -13'd86,  
13'd413,  -13'd38,  13'd1225,  -13'd316,  13'd1100,  -13'd351,  -13'd633,  -13'd398,  13'd392,  13'd436,  -13'd120,  13'd654,  13'd593,  13'd35,  -13'd281,  -13'd37,  
13'd825,  13'd380,  13'd228,  -13'd585,  -13'd1091,  13'd250,  13'd460,  -13'd530,  13'd78,  13'd352,  -13'd312,  13'd491,  -13'd182,  13'd427,  13'd302,  13'd496,  
13'd579,  -13'd485,  13'd871,  13'd732,  -13'd775,  -13'd495,  13'd284,  13'd339,  13'd52,  -13'd542,  13'd1030,  13'd794,  -13'd489,  -13'd345,  13'd231,  13'd277,  
-13'd420,  13'd129,  13'd516,  13'd693,  13'd813,  -13'd454,  13'd405,  -13'd631,  13'd869,  -13'd280,  -13'd216,  13'd301,  13'd141,  -13'd551,  -13'd455,  -13'd276,  
-13'd210,  13'd113,  -13'd1248,  13'd44,  13'd150,  -13'd300,  13'd137,  13'd572,  -13'd320,  13'd172,  13'd97,  13'd866,  13'd26,  -13'd230,  13'd219,  13'd293,  
13'd346,  13'd467,  -13'd457,  -13'd867,  -13'd1,  -13'd338,  -13'd78,  -13'd396,  13'd58,  13'd304,  -13'd751,  -13'd248,  13'd454,  13'd618,  13'd865,  13'd457,  
13'd646,  13'd287,  13'd924,  -13'd268,  13'd635,  -13'd60,  -13'd287,  -13'd21,  -13'd566,  13'd76,  -13'd707,  13'd25,  -13'd353,  13'd1126,  13'd147,  -13'd375,  
-13'd204,  13'd858,  -13'd14,  -13'd474,  -13'd848,  -13'd55,  13'd73,  -13'd158,  -13'd732,  -13'd41,  13'd601,  -13'd176,  -13'd78,  -13'd1080,  13'd726,  -13'd43,  
-13'd798,  13'd283,  -13'd333,  13'd367,  -13'd593,  -13'd214,  -13'd731,  13'd281,  13'd345,  -13'd494,  13'd494,  -13'd325,  13'd176,  13'd2,  13'd261,  -13'd549,  
13'd433,  13'd562,  -13'd3,  -13'd291,  -13'd68,  13'd436,  -13'd315,  -13'd677,  13'd375,  13'd257,  13'd70,  -13'd374,  -13'd187,  13'd74,  13'd538,  -13'd118,  
-13'd415,  13'd366,  -13'd494,  13'd842,  13'd565,  13'd674,  -13'd161,  13'd316,  13'd8,  13'd218,  13'd624,  13'd50,  13'd737,  -13'd251,  13'd147,  13'd146,  

-13'd620,  13'd700,  13'd236,  13'd137,  13'd449,  -13'd91,  -13'd1118,  13'd379,  13'd23,  13'd547,  13'd822,  -13'd238,  -13'd115,  -13'd375,  13'd414,  -13'd16,  
-13'd501,  -13'd477,  -13'd666,  13'd671,  13'd769,  -13'd102,  -13'd248,  13'd313,  13'd214,  13'd204,  13'd847,  -13'd54,  13'd646,  13'd641,  -13'd13,  13'd392,  
-13'd868,  13'd581,  13'd2,  13'd318,  13'd45,  13'd380,  -13'd87,  13'd347,  13'd110,  -13'd449,  -13'd6,  13'd238,  13'd365,  -13'd778,  13'd364,  13'd961,  
-13'd747,  -13'd274,  -13'd827,  13'd163,  -13'd195,  -13'd464,  -13'd572,  13'd267,  -13'd288,  13'd117,  -13'd99,  -13'd154,  13'd805,  -13'd402,  13'd368,  13'd402,  
13'd30,  -13'd758,  13'd431,  13'd86,  -13'd51,  13'd469,  13'd320,  -13'd60,  -13'd800,  -13'd394,  13'd344,  13'd137,  13'd386,  -13'd600,  -13'd758,  13'd362,  
-13'd94,  -13'd70,  13'd21,  13'd216,  13'd229,  13'd53,  -13'd32,  13'd651,  -13'd571,  13'd386,  -13'd43,  13'd464,  13'd104,  13'd79,  -13'd224,  13'd427,  
-13'd167,  -13'd728,  -13'd305,  13'd154,  -13'd463,  -13'd130,  13'd31,  13'd702,  -13'd786,  13'd14,  13'd627,  -13'd168,  13'd93,  -13'd449,  -13'd251,  -13'd203,  
-13'd524,  13'd175,  13'd209,  -13'd127,  -13'd52,  -13'd58,  -13'd147,  13'd138,  -13'd410,  13'd273,  13'd43,  -13'd350,  -13'd345,  13'd814,  -13'd546,  13'd642,  
-13'd232,  13'd881,  13'd410,  13'd354,  -13'd118,  -13'd276,  13'd631,  13'd256,  -13'd448,  -13'd104,  13'd40,  13'd716,  13'd319,  13'd342,  13'd239,  -13'd85,  
13'd21,  13'd773,  13'd253,  -13'd98,  13'd392,  -13'd245,  -13'd623,  13'd761,  -13'd802,  -13'd87,  -13'd154,  -13'd170,  -13'd477,  -13'd145,  13'd378,  13'd312,  
13'd203,  -13'd54,  -13'd285,  -13'd29,  -13'd850,  13'd121,  -13'd163,  -13'd833,  13'd626,  13'd130,  13'd249,  -13'd29,  -13'd622,  -13'd638,  -13'd760,  -13'd237,  
13'd455,  -13'd712,  -13'd185,  -13'd78,  -13'd184,  -13'd397,  13'd398,  13'd41,  -13'd10,  13'd98,  13'd487,  -13'd412,  13'd418,  -13'd277,  13'd45,  -13'd19,  
-13'd142,  -13'd378,  -13'd227,  13'd8,  -13'd34,  -13'd87,  13'd367,  -13'd81,  13'd468,  13'd323,  -13'd58,  -13'd323,  13'd355,  13'd491,  -13'd613,  13'd317,  
13'd768,  13'd380,  13'd448,  13'd155,  13'd295,  -13'd733,  13'd78,  13'd346,  -13'd40,  -13'd948,  -13'd444,  -13'd526,  -13'd711,  -13'd246,  13'd452,  -13'd544,  
-13'd253,  13'd205,  13'd547,  13'd249,  13'd972,  13'd403,  -13'd34,  -13'd93,  13'd434,  -13'd175,  -13'd577,  13'd374,  13'd519,  13'd298,  -13'd63,  -13'd267,  
-13'd204,  -13'd56,  -13'd414,  -13'd188,  13'd372,  13'd188,  13'd131,  13'd16,  13'd500,  13'd540,  13'd509,  13'd95,  13'd514,  -13'd539,  13'd84,  -13'd113,  
-13'd162,  -13'd322,  -13'd556,  13'd220,  -13'd171,  13'd278,  -13'd46,  -13'd2,  13'd501,  13'd452,  13'd73,  -13'd162,  13'd358,  13'd147,  13'd402,  -13'd361,  
13'd528,  13'd78,  -13'd136,  13'd330,  -13'd239,  13'd398,  -13'd264,  -13'd480,  13'd211,  13'd286,  -13'd234,  13'd60,  13'd366,  13'd1226,  -13'd183,  13'd315,  
-13'd365,  -13'd223,  13'd591,  13'd499,  13'd51,  -13'd152,  13'd141,  -13'd578,  13'd362,  -13'd340,  13'd79,  13'd690,  13'd174,  -13'd135,  -13'd184,  -13'd311,  
-13'd246,  -13'd594,  13'd107,  13'd288,  13'd845,  -13'd314,  -13'd222,  13'd110,  13'd267,  13'd592,  -13'd58,  13'd507,  13'd542,  13'd158,  13'd89,  -13'd530,  
13'd28,  -13'd85,  13'd95,  -13'd460,  -13'd944,  -13'd256,  13'd570,  13'd28,  13'd143,  -13'd272,  13'd799,  -13'd639,  -13'd354,  13'd427,  -13'd219,  -13'd64,  
13'd24,  13'd200,  -13'd282,  13'd594,  -13'd332,  13'd538,  13'd919,  13'd880,  13'd270,  13'd221,  13'd669,  -13'd236,  13'd84,  13'd502,  13'd982,  13'd39,  
-13'd203,  -13'd561,  13'd441,  13'd358,  -13'd458,  -13'd627,  -13'd387,  -13'd389,  -13'd556,  -13'd454,  -13'd705,  -13'd363,  -13'd492,  13'd1014,  13'd522,  13'd340,  
-13'd707,  13'd200,  -13'd208,  -13'd105,  13'd35,  -13'd142,  13'd302,  -13'd127,  -13'd36,  -13'd231,  -13'd125,  -13'd208,  13'd357,  -13'd295,  13'd268,  13'd331,  
13'd38,  13'd1102,  -13'd86,  13'd177,  13'd768,  13'd567,  -13'd606,  -13'd337,  13'd170,  13'd661,  13'd127,  -13'd105,  -13'd228,  13'd393,  -13'd598,  13'd175,  

-13'd761,  -13'd28,  -13'd101,  -13'd115,  -13'd428,  13'd318,  13'd701,  13'd349,  -13'd570,  13'd139,  13'd252,  13'd102,  13'd248,  13'd538,  13'd121,  -13'd425,  
13'd708,  -13'd88,  13'd44,  -13'd65,  13'd404,  13'd344,  13'd642,  13'd353,  -13'd440,  13'd300,  13'd1046,  13'd657,  -13'd133,  13'd232,  13'd202,  13'd227,  
13'd321,  13'd112,  -13'd79,  13'd582,  13'd754,  13'd264,  13'd443,  13'd76,  13'd264,  -13'd121,  13'd642,  13'd267,  -13'd76,  13'd523,  13'd483,  -13'd342,  
-13'd40,  13'd1130,  13'd721,  -13'd58,  -13'd148,  13'd95,  -13'd512,  13'd187,  13'd158,  -13'd244,  -13'd269,  13'd470,  13'd277,  -13'd474,  -13'd572,  13'd706,  
-13'd106,  13'd184,  13'd348,  -13'd145,  -13'd65,  13'd2,  -13'd861,  13'd197,  13'd474,  13'd312,  13'd33,  13'd30,  -13'd62,  13'd400,  -13'd389,  -13'd227,  
13'd273,  -13'd188,  -13'd650,  -13'd23,  -13'd39,  -13'd816,  13'd15,  13'd10,  -13'd528,  -13'd117,  13'd604,  -13'd446,  13'd9,  13'd146,  -13'd480,  -13'd96,  
-13'd395,  -13'd97,  13'd1011,  13'd433,  -13'd414,  13'd701,  13'd1101,  -13'd421,  13'd41,  13'd161,  -13'd315,  -13'd50,  -13'd709,  13'd141,  13'd203,  -13'd420,  
-13'd722,  13'd940,  13'd23,  13'd70,  13'd634,  -13'd52,  13'd526,  -13'd289,  13'd528,  13'd285,  13'd568,  -13'd1006,  -13'd174,  -13'd37,  -13'd285,  -13'd445,  
-13'd1152,  -13'd35,  -13'd479,  -13'd489,  13'd728,  -13'd306,  -13'd1024,  -13'd321,  -13'd141,  13'd781,  -13'd278,  -13'd336,  -13'd743,  -13'd395,  13'd127,  -13'd60,  
-13'd2070,  -13'd967,  13'd673,  -13'd648,  -13'd781,  13'd4,  -13'd623,  -13'd177,  -13'd423,  -13'd216,  -13'd36,  -13'd757,  -13'd986,  -13'd57,  13'd912,  13'd118,  
-13'd40,  -13'd563,  -13'd325,  -13'd285,  -13'd681,  -13'd419,  13'd1289,  -13'd448,  13'd331,  -13'd458,  -13'd41,  13'd332,  -13'd405,  -13'd310,  13'd15,  13'd228,  
13'd697,  -13'd606,  13'd92,  13'd60,  -13'd701,  -13'd404,  -13'd694,  13'd188,  13'd68,  13'd59,  -13'd488,  -13'd460,  -13'd133,  -13'd237,  -13'd732,  -13'd199,  
-13'd849,  -13'd57,  -13'd24,  -13'd113,  13'd266,  -13'd832,  -13'd596,  13'd228,  13'd526,  13'd476,  -13'd853,  -13'd140,  -13'd816,  13'd170,  -13'd70,  -13'd278,  
-13'd242,  13'd470,  13'd284,  -13'd70,  -13'd440,  13'd203,  13'd95,  -13'd1007,  13'd570,  -13'd449,  -13'd737,  13'd159,  -13'd429,  13'd593,  -13'd245,  -13'd913,  
-13'd317,  -13'd143,  13'd1025,  13'd64,  -13'd296,  -13'd117,  -13'd79,  -13'd68,  13'd548,  13'd65,  -13'd771,  13'd1198,  -13'd751,  13'd623,  13'd494,  -13'd1117,  
13'd858,  13'd355,  13'd393,  -13'd177,  -13'd812,  13'd258,  13'd23,  13'd358,  13'd44,  13'd655,  -13'd813,  13'd51,  13'd742,  13'd352,  13'd199,  13'd64,  
-13'd166,  -13'd9,  13'd228,  -13'd298,  -13'd600,  13'd449,  13'd285,  13'd500,  13'd357,  -13'd120,  13'd460,  13'd405,  -13'd385,  13'd1161,  13'd581,  13'd906,  
13'd232,  -13'd793,  13'd275,  13'd391,  -13'd364,  13'd300,  -13'd178,  13'd268,  -13'd236,  13'd126,  13'd172,  13'd328,  13'd55,  13'd261,  -13'd252,  13'd686,  
13'd49,  13'd401,  13'd576,  13'd614,  -13'd168,  -13'd51,  13'd156,  -13'd409,  13'd173,  -13'd272,  -13'd93,  13'd50,  13'd535,  13'd387,  13'd264,  -13'd264,  
13'd1339,  -13'd5,  13'd487,  13'd809,  13'd309,  -13'd301,  13'd165,  -13'd47,  -13'd607,  13'd502,  13'd326,  13'd712,  13'd766,  -13'd747,  13'd80,  -13'd604,  
-13'd135,  -13'd123,  -13'd304,  13'd191,  -13'd298,  -13'd431,  -13'd23,  -13'd227,  -13'd511,  -13'd106,  -13'd411,  -13'd56,  -13'd218,  13'd34,  -13'd63,  13'd186,  
-13'd434,  13'd336,  -13'd175,  13'd596,  13'd10,  13'd62,  13'd424,  -13'd619,  -13'd173,  13'd68,  13'd166,  -13'd185,  -13'd86,  13'd825,  13'd417,  13'd76,  
-13'd37,  13'd478,  13'd471,  13'd208,  -13'd149,  13'd221,  13'd415,  13'd236,  13'd242,  13'd218,  -13'd11,  -13'd308,  -13'd155,  -13'd481,  -13'd358,  13'd109,  
-13'd147,  13'd807,  -13'd288,  -13'd165,  13'd33,  -13'd320,  -13'd502,  13'd119,  13'd64,  -13'd632,  -13'd1,  -13'd834,  13'd417,  -13'd472,  -13'd155,  13'd719,  
-13'd237,  13'd474,  -13'd868,  -13'd153,  13'd355,  -13'd318,  -13'd123,  13'd340,  -13'd449,  13'd20,  -13'd390,  -13'd162,  -13'd137,  -13'd131,  -13'd210,  13'd62,  

-13'd144,  13'd756,  -13'd256,  -13'd157,  13'd119,  -13'd53,  -13'd339,  -13'd101,  13'd274,  13'd113,  -13'd325,  -13'd166,  13'd713,  -13'd603,  13'd185,  13'd281,  
-13'd275,  -13'd183,  -13'd763,  13'd94,  13'd226,  13'd466,  -13'd495,  13'd138,  -13'd132,  -13'd353,  -13'd626,  13'd184,  13'd518,  -13'd169,  13'd571,  13'd446,  
-13'd272,  -13'd398,  13'd315,  13'd278,  -13'd276,  -13'd278,  13'd660,  13'd56,  -13'd731,  -13'd25,  13'd418,  -13'd162,  13'd355,  -13'd1021,  13'd51,  13'd194,  
-13'd384,  -13'd294,  -13'd290,  -13'd216,  -13'd303,  13'd365,  13'd772,  -13'd558,  13'd378,  -13'd32,  13'd584,  13'd347,  -13'd714,  13'd471,  -13'd476,  13'd199,  
-13'd189,  13'd531,  -13'd480,  13'd24,  -13'd319,  -13'd242,  13'd518,  13'd20,  -13'd332,  -13'd412,  13'd18,  -13'd41,  -13'd590,  13'd65,  -13'd835,  13'd54,  
13'd214,  13'd101,  13'd24,  13'd693,  -13'd49,  -13'd179,  -13'd557,  13'd612,  -13'd436,  -13'd1146,  13'd419,  13'd99,  -13'd374,  13'd370,  -13'd110,  13'd336,  
-13'd568,  13'd253,  13'd15,  -13'd164,  13'd121,  13'd588,  -13'd138,  -13'd66,  -13'd498,  13'd193,  13'd530,  -13'd59,  13'd526,  -13'd870,  13'd531,  13'd645,  
-13'd185,  13'd2,  -13'd673,  -13'd544,  13'd761,  -13'd486,  13'd148,  -13'd109,  13'd212,  -13'd265,  13'd601,  13'd56,  -13'd343,  -13'd424,  -13'd57,  13'd800,  
13'd132,  -13'd219,  -13'd333,  -13'd488,  -13'd303,  13'd344,  13'd496,  13'd184,  13'd436,  13'd430,  13'd131,  -13'd323,  -13'd30,  13'd296,  -13'd144,  -13'd262,  
13'd523,  13'd686,  13'd629,  13'd449,  13'd17,  -13'd300,  -13'd522,  13'd305,  -13'd52,  13'd652,  13'd78,  -13'd748,  13'd567,  13'd268,  -13'd183,  -13'd268,  
13'd485,  13'd18,  13'd332,  -13'd364,  -13'd687,  -13'd391,  -13'd486,  13'd271,  13'd313,  13'd117,  13'd378,  -13'd663,  13'd642,  13'd208,  13'd66,  -13'd212,  
-13'd174,  13'd336,  -13'd212,  13'd21,  13'd431,  -13'd64,  -13'd861,  -13'd23,  -13'd498,  13'd145,  13'd75,  13'd415,  13'd314,  -13'd384,  -13'd343,  13'd140,  
-13'd633,  -13'd437,  13'd687,  -13'd388,  -13'd83,  13'd581,  -13'd389,  -13'd53,  -13'd753,  -13'd154,  -13'd269,  13'd39,  13'd459,  -13'd25,  13'd466,  -13'd422,  
-13'd327,  -13'd489,  -13'd695,  13'd313,  13'd392,  13'd146,  13'd4,  -13'd806,  13'd83,  13'd486,  -13'd214,  -13'd283,  13'd212,  -13'd840,  13'd31,  13'd271,  
-13'd959,  -13'd460,  13'd469,  13'd402,  -13'd59,  -13'd26,  -13'd602,  -13'd4,  13'd418,  13'd1162,  -13'd7,  13'd312,  -13'd489,  13'd679,  -13'd482,  -13'd480,  
-13'd896,  13'd203,  -13'd47,  13'd19,  -13'd98,  -13'd22,  -13'd434,  -13'd246,  13'd1209,  -13'd32,  13'd496,  -13'd1022,  -13'd496,  -13'd797,  -13'd415,  -13'd832,  
-13'd511,  -13'd271,  -13'd584,  -13'd320,  -13'd504,  13'd185,  -13'd418,  -13'd337,  -13'd258,  13'd824,  13'd668,  -13'd640,  13'd234,  -13'd659,  -13'd625,  -13'd446,  
-13'd44,  -13'd148,  13'd334,  -13'd161,  13'd187,  -13'd322,  -13'd247,  -13'd45,  -13'd277,  -13'd132,  13'd78,  -13'd163,  -13'd270,  -13'd553,  -13'd186,  13'd328,  
-13'd233,  -13'd6,  -13'd426,  13'd472,  13'd792,  13'd500,  -13'd681,  13'd55,  -13'd373,  -13'd526,  -13'd346,  13'd522,  13'd789,  -13'd555,  -13'd131,  13'd182,  
-13'd712,  -13'd135,  13'd144,  13'd598,  -13'd76,  13'd344,  13'd238,  -13'd226,  13'd334,  13'd428,  -13'd102,  13'd278,  13'd81,  13'd169,  -13'd504,  -13'd606,  
-13'd148,  -13'd181,  -13'd620,  13'd510,  13'd214,  13'd340,  13'd1129,  -13'd440,  13'd607,  13'd189,  13'd885,  -13'd430,  -13'd229,  -13'd307,  -13'd65,  -13'd508,  
13'd623,  13'd84,  -13'd128,  -13'd96,  -13'd470,  -13'd659,  13'd34,  -13'd571,  13'd1112,  13'd795,  -13'd88,  13'd442,  13'd324,  -13'd1140,  -13'd220,  13'd39,  
13'd285,  13'd555,  -13'd341,  13'd450,  13'd6,  13'd38,  -13'd254,  -13'd56,  13'd766,  13'd1002,  13'd434,  13'd615,  -13'd354,  13'd180,  -13'd402,  13'd530,  
13'd805,  13'd551,  -13'd523,  -13'd425,  13'd503,  13'd602,  -13'd236,  13'd381,  13'd350,  -13'd419,  -13'd53,  -13'd450,  13'd761,  13'd649,  -13'd121,  -13'd300,  
13'd201,  13'd162,  13'd748,  13'd203,  -13'd97,  13'd371,  -13'd309,  -13'd479,  13'd713,  13'd124,  -13'd190,  -13'd492,  -13'd109,  13'd531,  -13'd570,  13'd361,  

13'd872,  -13'd876,  -13'd485,  13'd56,  -13'd765,  13'd442,  13'd192,  -13'd273,  -13'd515,  13'd293,  13'd621,  13'd107,  -13'd379,  13'd422,  -13'd792,  -13'd370,  
-13'd203,  -13'd343,  -13'd64,  -13'd651,  -13'd556,  13'd178,  13'd125,  -13'd1052,  13'd60,  -13'd120,  -13'd139,  13'd762,  -13'd160,  13'd251,  13'd165,  13'd71,  
13'd349,  13'd1,  -13'd86,  -13'd284,  13'd330,  -13'd266,  -13'd657,  13'd583,  13'd716,  -13'd150,  -13'd187,  13'd367,  13'd279,  -13'd186,  -13'd151,  13'd619,  
-13'd42,  13'd169,  -13'd208,  13'd260,  -13'd263,  -13'd82,  13'd158,  13'd220,  13'd369,  -13'd368,  -13'd770,  -13'd362,  -13'd598,  13'd248,  13'd329,  13'd379,  
-13'd585,  13'd162,  -13'd1,  13'd83,  13'd85,  -13'd134,  13'd539,  13'd25,  13'd286,  -13'd55,  -13'd621,  13'd179,  13'd1,  13'd359,  -13'd651,  -13'd460,  
13'd102,  -13'd152,  13'd212,  13'd349,  13'd191,  13'd390,  13'd878,  -13'd468,  13'd748,  -13'd295,  13'd201,  13'd721,  -13'd42,  13'd385,  -13'd468,  -13'd556,  
13'd131,  13'd283,  13'd160,  13'd335,  -13'd6,  -13'd104,  13'd469,  -13'd577,  13'd986,  13'd422,  -13'd959,  13'd120,  -13'd156,  13'd522,  13'd641,  13'd566,  
13'd682,  13'd566,  13'd76,  -13'd24,  13'd512,  -13'd131,  13'd631,  13'd90,  -13'd536,  -13'd291,  -13'd198,  13'd320,  -13'd355,  -13'd124,  13'd182,  -13'd6,  
-13'd484,  -13'd390,  13'd24,  13'd71,  13'd518,  -13'd325,  13'd13,  -13'd754,  13'd398,  -13'd237,  -13'd775,  13'd436,  -13'd10,  13'd382,  -13'd438,  13'd419,  
13'd817,  -13'd236,  -13'd677,  13'd644,  -13'd320,  -13'd659,  13'd543,  -13'd300,  13'd8,  -13'd725,  13'd370,  13'd255,  13'd233,  -13'd72,  13'd287,  13'd423,  
13'd369,  13'd223,  13'd1004,  13'd86,  13'd260,  13'd156,  13'd517,  13'd413,  -13'd396,  13'd207,  -13'd957,  13'd748,  13'd156,  13'd268,  13'd70,  13'd618,  
13'd310,  13'd101,  13'd88,  13'd96,  13'd743,  -13'd55,  13'd110,  13'd373,  13'd202,  13'd153,  -13'd420,  13'd206,  13'd175,  13'd123,  -13'd498,  -13'd126,  
13'd352,  -13'd64,  -13'd145,  13'd237,  -13'd874,  13'd489,  13'd493,  13'd87,  -13'd553,  -13'd724,  -13'd321,  13'd215,  -13'd804,  -13'd365,  -13'd303,  13'd322,  
13'd363,  -13'd60,  -13'd578,  -13'd52,  -13'd636,  13'd363,  13'd43,  13'd56,  13'd113,  -13'd245,  13'd3,  13'd186,  13'd381,  13'd494,  -13'd184,  -13'd345,  
-13'd5,  -13'd8,  -13'd534,  -13'd4,  13'd606,  13'd467,  -13'd25,  -13'd308,  -13'd582,  -13'd188,  13'd31,  -13'd213,  13'd881,  -13'd26,  -13'd417,  13'd405,  
13'd473,  13'd229,  13'd695,  13'd62,  13'd388,  -13'd31,  13'd144,  13'd341,  -13'd634,  13'd390,  -13'd956,  13'd811,  13'd494,  13'd325,  13'd340,  13'd7,  
13'd349,  13'd601,  -13'd21,  -13'd612,  -13'd162,  13'd32,  13'd123,  -13'd0,  -13'd545,  13'd85,  -13'd481,  -13'd764,  13'd681,  13'd145,  -13'd107,  13'd467,  
13'd717,  -13'd21,  -13'd347,  -13'd233,  -13'd457,  -13'd516,  13'd54,  13'd577,  -13'd344,  -13'd226,  13'd16,  -13'd454,  -13'd722,  13'd360,  -13'd265,  13'd232,  
13'd35,  13'd51,  -13'd203,  -13'd460,  13'd616,  -13'd916,  13'd608,  -13'd78,  -13'd386,  -13'd31,  13'd55,  -13'd294,  -13'd627,  -13'd691,  13'd150,  13'd345,  
-13'd674,  -13'd460,  -13'd206,  13'd629,  -13'd244,  -13'd449,  -13'd246,  -13'd400,  13'd77,  -13'd306,  13'd313,  13'd79,  -13'd677,  -13'd160,  -13'd387,  13'd131,  
13'd509,  13'd82,  13'd97,  13'd660,  -13'd307,  13'd518,  -13'd518,  13'd171,  -13'd1323,  13'd736,  -13'd532,  -13'd54,  -13'd282,  13'd1011,  13'd111,  -13'd76,  
13'd269,  -13'd538,  13'd433,  -13'd179,  -13'd653,  -13'd523,  -13'd401,  13'd611,  13'd54,  13'd42,  -13'd502,  -13'd265,  13'd307,  13'd676,  -13'd392,  -13'd131,  
-13'd330,  13'd196,  13'd8,  13'd253,  -13'd8,  13'd90,  -13'd875,  13'd490,  -13'd243,  -13'd466,  -13'd548,  -13'd291,  13'd432,  13'd214,  13'd728,  -13'd405,  
13'd52,  -13'd327,  13'd324,  13'd301,  13'd553,  -13'd436,  -13'd268,  -13'd232,  -13'd817,  -13'd487,  13'd63,  -13'd498,  -13'd401,  -13'd545,  13'd497,  -13'd331,  
-13'd209,  -13'd200,  -13'd246,  13'd108,  13'd129,  13'd544,  13'd139,  13'd179,  -13'd535,  -13'd961,  13'd140,  13'd431,  -13'd85,  -13'd182,  13'd542,  -13'd215,  

-13'd732,  -13'd423,  13'd68,  -13'd311,  -13'd723,  -13'd218,  13'd558,  13'd272,  13'd413,  -13'd186,  -13'd650,  -13'd271,  -13'd1061,  -13'd47,  -13'd247,  -13'd951,  
-13'd511,  13'd119,  -13'd817,  13'd523,  13'd37,  -13'd34,  13'd83,  13'd226,  13'd527,  -13'd440,  -13'd233,  -13'd360,  -13'd386,  -13'd32,  13'd469,  -13'd277,  
13'd172,  -13'd490,  13'd328,  -13'd415,  -13'd407,  -13'd199,  -13'd1011,  -13'd225,  13'd470,  13'd75,  -13'd212,  -13'd233,  13'd113,  -13'd438,  -13'd334,  13'd91,  
-13'd633,  -13'd86,  -13'd239,  13'd155,  13'd378,  -13'd740,  -13'd241,  13'd577,  -13'd703,  13'd490,  -13'd532,  13'd13,  13'd766,  -13'd1097,  13'd96,  13'd650,  
-13'd561,  -13'd1092,  13'd312,  -13'd142,  13'd548,  13'd105,  -13'd22,  -13'd124,  13'd138,  -13'd701,  13'd20,  -13'd258,  -13'd21,  13'd716,  13'd487,  13'd134,  
-13'd213,  -13'd380,  -13'd782,  -13'd168,  13'd172,  -13'd477,  13'd163,  -13'd32,  -13'd83,  -13'd144,  -13'd139,  -13'd190,  -13'd277,  13'd10,  -13'd919,  -13'd478,  
-13'd236,  13'd101,  -13'd143,  -13'd341,  -13'd44,  -13'd430,  -13'd1098,  -13'd307,  -13'd639,  13'd911,  13'd11,  13'd330,  -13'd668,  13'd335,  -13'd774,  13'd732,  
-13'd124,  -13'd224,  -13'd386,  -13'd637,  13'd335,  13'd519,  -13'd186,  13'd481,  13'd551,  13'd298,  -13'd408,  13'd793,  13'd112,  13'd26,  13'd705,  -13'd483,  
-13'd437,  -13'd951,  -13'd553,  13'd195,  -13'd373,  13'd388,  -13'd322,  -13'd115,  -13'd237,  -13'd244,  13'd166,  13'd24,  -13'd150,  -13'd515,  13'd67,  13'd481,  
-13'd95,  -13'd99,  13'd544,  13'd460,  13'd373,  13'd317,  13'd363,  13'd530,  -13'd704,  -13'd183,  13'd725,  13'd743,  13'd918,  -13'd575,  -13'd20,  13'd465,  
13'd263,  13'd102,  -13'd555,  13'd566,  13'd105,  13'd424,  -13'd52,  13'd111,  13'd525,  -13'd647,  -13'd1234,  13'd34,  13'd462,  -13'd468,  -13'd82,  -13'd548,  
-13'd656,  13'd381,  13'd511,  -13'd500,  -13'd190,  13'd334,  13'd248,  -13'd678,  13'd462,  13'd180,  13'd150,  13'd272,  -13'd147,  -13'd365,  13'd434,  -13'd662,  
13'd277,  13'd204,  13'd360,  -13'd391,  13'd46,  -13'd248,  -13'd318,  -13'd954,  -13'd496,  13'd898,  13'd784,  13'd354,  -13'd40,  13'd7,  -13'd50,  13'd289,  
13'd400,  13'd41,  13'd509,  13'd38,  -13'd125,  -13'd562,  13'd182,  13'd740,  -13'd39,  13'd305,  13'd436,  -13'd371,  -13'd21,  13'd758,  -13'd592,  13'd416,  
-13'd192,  -13'd352,  -13'd1036,  -13'd503,  13'd419,  -13'd238,  -13'd231,  -13'd4,  -13'd835,  -13'd179,  13'd88,  -13'd670,  13'd244,  13'd182,  13'd490,  13'd656,  
13'd530,  -13'd131,  13'd298,  13'd375,  13'd383,  13'd805,  -13'd625,  -13'd228,  13'd878,  -13'd112,  -13'd327,  -13'd398,  -13'd594,  -13'd80,  13'd465,  -13'd375,  
-13'd468,  13'd424,  13'd288,  -13'd7,  13'd192,  13'd343,  -13'd545,  -13'd462,  13'd932,  13'd319,  13'd220,  -13'd720,  -13'd328,  -13'd355,  -13'd24,  13'd145,  
13'd504,  -13'd233,  -13'd121,  13'd237,  13'd830,  -13'd37,  13'd236,  13'd417,  -13'd123,  -13'd300,  13'd61,  13'd264,  -13'd138,  -13'd19,  13'd37,  13'd411,  
-13'd431,  -13'd156,  -13'd256,  -13'd354,  13'd315,  -13'd557,  13'd712,  -13'd684,  13'd340,  13'd383,  -13'd27,  13'd147,  -13'd95,  13'd65,  13'd176,  -13'd354,  
-13'd442,  -13'd865,  -13'd120,  -13'd458,  -13'd920,  -13'd135,  -13'd440,  -13'd74,  -13'd809,  -13'd987,  -13'd621,  -13'd105,  -13'd768,  13'd102,  -13'd499,  -13'd497,  
-13'd170,  -13'd229,  13'd320,  13'd313,  13'd998,  13'd336,  -13'd129,  13'd335,  13'd173,  -13'd346,  13'd523,  -13'd183,  13'd636,  -13'd157,  -13'd110,  -13'd448,  
13'd29,  13'd15,  13'd350,  13'd129,  13'd571,  -13'd132,  -13'd561,  13'd83,  -13'd692,  -13'd465,  13'd31,  -13'd185,  13'd142,  -13'd993,  13'd318,  -13'd288,  
13'd397,  -13'd383,  13'd436,  13'd320,  -13'd884,  13'd639,  13'd376,  -13'd526,  -13'd288,  -13'd927,  13'd258,  -13'd18,  -13'd155,  -13'd197,  -13'd372,  -13'd260,  
-13'd53,  -13'd462,  13'd51,  13'd695,  -13'd657,  13'd693,  13'd566,  -13'd893,  13'd849,  -13'd1237,  -13'd313,  13'd601,  -13'd881,  13'd205,  -13'd555,  -13'd360,  
13'd167,  -13'd188,  13'd1610,  13'd132,  -13'd427,  13'd39,  -13'd39,  -13'd469,  13'd1417,  13'd739,  -13'd43,  -13'd608,  -13'd666,  13'd606,  -13'd1335,  -13'd664,  

13'd74,  13'd243,  -13'd670,  13'd288,  -13'd536,  13'd89,  13'd648,  13'd276,  13'd287,  13'd172,  -13'd356,  -13'd314,  13'd54,  13'd347,  13'd58,  13'd324,  
13'd376,  -13'd416,  -13'd359,  -13'd283,  -13'd64,  13'd11,  13'd547,  -13'd495,  13'd889,  13'd248,  -13'd767,  -13'd215,  13'd164,  13'd526,  13'd813,  -13'd34,  
-13'd475,  -13'd66,  13'd7,  -13'd572,  13'd36,  -13'd437,  13'd421,  -13'd289,  -13'd562,  13'd355,  13'd77,  13'd299,  -13'd230,  -13'd94,  -13'd481,  13'd343,  
-13'd254,  13'd377,  13'd280,  -13'd54,  -13'd186,  -13'd769,  13'd428,  -13'd278,  13'd416,  -13'd662,  13'd126,  13'd287,  13'd239,  -13'd13,  -13'd427,  13'd746,  
13'd227,  13'd1038,  -13'd456,  13'd580,  13'd577,  13'd36,  13'd58,  13'd416,  -13'd376,  13'd103,  13'd134,  13'd88,  13'd103,  -13'd341,  13'd448,  13'd588,  
-13'd456,  13'd639,  13'd144,  13'd98,  13'd9,  -13'd466,  13'd444,  13'd195,  -13'd218,  13'd710,  -13'd208,  -13'd815,  13'd331,  13'd337,  13'd452,  -13'd185,  
-13'd217,  -13'd825,  -13'd14,  13'd183,  13'd441,  13'd159,  -13'd686,  13'd32,  -13'd1117,  13'd654,  -13'd276,  -13'd308,  13'd227,  13'd1208,  13'd579,  -13'd377,  
13'd194,  -13'd329,  -13'd27,  13'd686,  13'd322,  -13'd158,  13'd531,  13'd892,  -13'd420,  -13'd754,  -13'd332,  13'd501,  -13'd127,  -13'd318,  13'd628,  13'd274,  
13'd45,  -13'd480,  13'd313,  13'd23,  -13'd208,  13'd24,  13'd543,  13'd539,  13'd691,  -13'd959,  13'd718,  13'd235,  -13'd115,  -13'd760,  13'd0,  -13'd725,  
13'd1107,  -13'd510,  -13'd950,  -13'd559,  13'd184,  13'd543,  13'd189,  13'd494,  -13'd366,  -13'd604,  13'd214,  -13'd732,  13'd451,  13'd145,  -13'd1169,  13'd191,  
-13'd615,  13'd289,  -13'd1021,  13'd430,  13'd836,  -13'd145,  -13'd424,  -13'd114,  -13'd34,  -13'd628,  -13'd462,  -13'd458,  13'd673,  -13'd782,  -13'd505,  -13'd588,  
-13'd350,  13'd633,  -13'd216,  13'd478,  13'd80,  13'd210,  -13'd896,  13'd237,  -13'd172,  13'd227,  -13'd49,  -13'd104,  -13'd381,  13'd794,  13'd383,  13'd429,  
13'd902,  13'd740,  -13'd285,  13'd310,  13'd240,  13'd343,  -13'd236,  -13'd21,  13'd64,  13'd596,  13'd255,  -13'd437,  13'd529,  -13'd704,  13'd209,  -13'd262,  
-13'd1114,  -13'd847,  -13'd575,  -13'd750,  13'd45,  -13'd766,  -13'd66,  -13'd38,  -13'd12,  -13'd150,  -13'd782,  -13'd966,  13'd514,  -13'd485,  -13'd387,  13'd51,  
-13'd782,  -13'd333,  -13'd643,  -13'd230,  -13'd77,  13'd26,  -13'd566,  13'd223,  -13'd624,  13'd414,  13'd450,  -13'd80,  -13'd605,  13'd86,  -13'd279,  13'd810,  
-13'd430,  -13'd498,  -13'd566,  13'd328,  13'd192,  -13'd167,  -13'd681,  -13'd675,  13'd143,  13'd379,  -13'd1005,  13'd337,  -13'd139,  13'd239,  -13'd25,  13'd328,  
13'd390,  13'd674,  13'd863,  13'd189,  13'd833,  -13'd212,  13'd495,  -13'd196,  -13'd397,  13'd529,  -13'd498,  -13'd35,  -13'd47,  13'd346,  -13'd425,  13'd102,  
13'd310,  13'd511,  13'd353,  -13'd334,  13'd288,  13'd129,  13'd53,  -13'd618,  -13'd769,  -13'd47,  -13'd862,  13'd442,  13'd239,  -13'd825,  13'd92,  13'd217,  
13'd55,  -13'd601,  -13'd362,  13'd41,  13'd726,  13'd520,  13'd100,  -13'd341,  13'd325,  -13'd205,  -13'd525,  13'd575,  13'd98,  13'd556,  -13'd365,  -13'd270,  
-13'd315,  -13'd5,  13'd1371,  -13'd395,  -13'd674,  -13'd10,  -13'd212,  -13'd151,  13'd82,  -13'd836,  -13'd170,  13'd310,  13'd19,  13'd530,  -13'd1173,  -13'd701,  
-13'd162,  -13'd121,  13'd90,  -13'd24,  13'd683,  -13'd20,  -13'd1127,  13'd239,  13'd1243,  -13'd548,  -13'd99,  -13'd92,  -13'd18,  -13'd1090,  13'd19,  -13'd94,  
13'd50,  -13'd204,  -13'd230,  13'd325,  13'd589,  13'd368,  -13'd371,  -13'd6,  13'd319,  13'd9,  13'd388,  13'd294,  13'd119,  -13'd1012,  -13'd609,  13'd528,  
13'd673,  13'd379,  -13'd13,  -13'd363,  13'd282,  13'd81,  -13'd340,  -13'd9,  13'd25,  13'd794,  13'd424,  13'd965,  13'd614,  -13'd496,  -13'd592,  -13'd638,  
13'd157,  13'd193,  13'd573,  -13'd117,  -13'd449,  13'd773,  13'd552,  13'd192,  13'd772,  13'd404,  13'd580,  13'd798,  13'd464,  13'd728,  -13'd275,  -13'd278,  
13'd94,  13'd153,  13'd258,  -13'd607,  13'd116,  13'd426,  13'd515,  13'd504,  13'd1184,  -13'd1196,  13'd160,  13'd322,  13'd542,  13'd964,  -13'd807,  -13'd18,  

-13'd372,  13'd87,  -13'd646,  -13'd793,  -13'd658,  -13'd436,  13'd333,  -13'd210,  -13'd206,  -13'd370,  13'd191,  -13'd20,  -13'd312,  -13'd585,  -13'd360,  -13'd35,  
-13'd172,  13'd638,  13'd169,  -13'd143,  -13'd412,  -13'd316,  -13'd155,  -13'd141,  13'd293,  13'd131,  -13'd333,  -13'd536,  13'd3,  13'd339,  13'd350,  13'd96,  
-13'd288,  13'd577,  13'd439,  13'd247,  -13'd568,  13'd297,  13'd351,  13'd529,  -13'd616,  13'd401,  -13'd505,  -13'd560,  13'd241,  -13'd946,  -13'd238,  13'd439,  
-13'd408,  -13'd627,  13'd479,  13'd114,  13'd253,  13'd293,  -13'd341,  13'd86,  -13'd510,  -13'd149,  -13'd336,  13'd5,  -13'd239,  13'd375,  13'd176,  -13'd55,  
-13'd542,  -13'd13,  -13'd538,  -13'd89,  -13'd253,  -13'd293,  13'd11,  -13'd51,  13'd132,  13'd273,  13'd369,  -13'd691,  -13'd654,  13'd453,  -13'd288,  -13'd311,  
-13'd529,  13'd513,  13'd327,  13'd214,  -13'd560,  -13'd445,  13'd113,  -13'd331,  -13'd99,  -13'd1110,  13'd820,  13'd484,  -13'd515,  13'd244,  13'd383,  -13'd612,  
13'd995,  13'd477,  13'd468,  13'd473,  -13'd186,  -13'd427,  13'd437,  13'd101,  13'd267,  -13'd402,  -13'd765,  -13'd52,  -13'd241,  13'd300,  13'd214,  -13'd476,  
13'd237,  -13'd356,  -13'd157,  -13'd216,  13'd101,  -13'd425,  -13'd378,  13'd268,  -13'd255,  -13'd381,  -13'd490,  13'd23,  13'd25,  -13'd731,  13'd223,  -13'd144,  
13'd301,  13'd100,  13'd10,  13'd252,  -13'd204,  -13'd439,  13'd87,  -13'd269,  -13'd586,  -13'd440,  -13'd91,  -13'd205,  -13'd295,  13'd306,  13'd366,  13'd682,  
-13'd321,  13'd822,  13'd861,  -13'd47,  -13'd344,  13'd82,  13'd176,  13'd911,  -13'd174,  13'd60,  -13'd446,  13'd40,  13'd178,  13'd213,  -13'd586,  13'd362,  
13'd415,  13'd72,  13'd397,  -13'd474,  -13'd788,  -13'd783,  13'd1104,  -13'd223,  13'd497,  -13'd129,  -13'd1149,  -13'd17,  13'd92,  13'd988,  13'd213,  -13'd590,  
13'd159,  13'd461,  13'd310,  -13'd30,  13'd138,  -13'd540,  13'd145,  13'd647,  13'd427,  13'd301,  -13'd651,  -13'd265,  -13'd610,  13'd282,  -13'd209,  13'd364,  
13'd145,  13'd705,  13'd91,  -13'd421,  -13'd371,  13'd393,  -13'd764,  13'd372,  -13'd355,  -13'd175,  -13'd600,  -13'd894,  13'd303,  13'd290,  13'd194,  -13'd117,  
13'd310,  13'd1006,  -13'd19,  -13'd84,  13'd742,  13'd101,  13'd127,  13'd14,  -13'd601,  13'd542,  13'd694,  -13'd33,  13'd217,  13'd491,  13'd441,  13'd114,  
13'd554,  -13'd326,  13'd633,  13'd598,  13'd601,  13'd583,  13'd355,  13'd741,  -13'd393,  -13'd496,  13'd219,  -13'd360,  13'd128,  -13'd296,  13'd232,  13'd292,  
-13'd974,  -13'd139,  13'd347,  13'd585,  13'd136,  13'd704,  13'd9,  13'd317,  -13'd1036,  -13'd230,  -13'd286,  -13'd268,  -13'd159,  13'd498,  -13'd405,  -13'd455,  
-13'd541,  13'd209,  13'd282,  13'd326,  13'd218,  -13'd321,  -13'd770,  13'd241,  -13'd1919,  13'd38,  13'd410,  -13'd210,  13'd33,  -13'd238,  -13'd165,  -13'd828,  
13'd112,  13'd311,  13'd118,  13'd211,  -13'd578,  -13'd64,  13'd17,  -13'd26,  -13'd1129,  -13'd185,  13'd568,  13'd190,  -13'd678,  -13'd767,  13'd242,  -13'd452,  
-13'd218,  13'd71,  -13'd320,  -13'd186,  -13'd538,  13'd456,  13'd448,  13'd322,  13'd246,  -13'd852,  13'd610,  13'd621,  13'd287,  -13'd310,  -13'd146,  13'd85,  
-13'd223,  -13'd191,  13'd129,  -13'd251,  -13'd173,  13'd282,  13'd721,  13'd652,  13'd9,  -13'd1099,  -13'd256,  -13'd649,  -13'd183,  13'd66,  -13'd371,  -13'd85,  
-13'd460,  13'd705,  -13'd193,  13'd484,  13'd681,  13'd346,  -13'd687,  13'd213,  13'd289,  13'd21,  13'd574,  -13'd77,  13'd38,  -13'd714,  -13'd97,  -13'd69,  
-13'd672,  13'd510,  -13'd197,  13'd693,  13'd488,  13'd81,  13'd524,  13'd328,  13'd819,  -13'd271,  13'd353,  -13'd4,  -13'd421,  -13'd775,  13'd19,  -13'd173,  
13'd361,  13'd23,  -13'd259,  13'd684,  13'd393,  -13'd409,  13'd826,  13'd255,  13'd860,  -13'd32,  -13'd170,  13'd40,  -13'd70,  -13'd81,  -13'd346,  -13'd361,  
13'd78,  -13'd36,  -13'd62,  13'd118,  -13'd78,  -13'd258,  -13'd292,  13'd309,  13'd338,  13'd598,  -13'd630,  13'd43,  13'd495,  13'd526,  13'd189,  -13'd484,  
-13'd231,  13'd48,  -13'd724,  -13'd1244,  -13'd473,  13'd167,  -13'd647,  -13'd727,  -13'd197,  -13'd392,  13'd166,  -13'd245,  -13'd442,  13'd405,  -13'd773,  -13'd116,  

-13'd51,  13'd547,  -13'd785,  -13'd323,  -13'd560,  13'd184,  -13'd160,  -13'd81,  -13'd162,  13'd33,  13'd536,  -13'd401,  -13'd492,  -13'd171,  13'd75,  13'd183,  
13'd137,  13'd168,  -13'd123,  13'd46,  -13'd431,  13'd824,  13'd466,  -13'd466,  -13'd133,  -13'd675,  -13'd204,  13'd84,  -13'd583,  13'd73,  -13'd907,  13'd295,  
-13'd606,  -13'd644,  -13'd625,  -13'd481,  13'd430,  13'd125,  13'd269,  13'd365,  13'd263,  13'd456,  13'd229,  13'd601,  13'd17,  13'd193,  13'd643,  -13'd394,  
13'd186,  13'd225,  13'd434,  -13'd596,  -13'd344,  -13'd488,  -13'd169,  13'd328,  13'd627,  13'd339,  -13'd28,  -13'd18,  -13'd231,  13'd772,  -13'd225,  13'd327,  
-13'd184,  13'd550,  13'd167,  13'd393,  13'd373,  13'd103,  13'd643,  -13'd291,  13'd362,  13'd589,  13'd430,  13'd413,  -13'd293,  -13'd232,  -13'd9,  -13'd756,  
13'd290,  -13'd86,  13'd137,  13'd350,  -13'd463,  13'd95,  13'd441,  -13'd45,  13'd735,  13'd904,  -13'd141,  13'd388,  -13'd188,  -13'd46,  -13'd351,  -13'd624,  
13'd84,  13'd258,  13'd277,  -13'd457,  13'd28,  13'd451,  13'd846,  13'd96,  13'd527,  -13'd471,  -13'd50,  13'd245,  -13'd211,  13'd823,  -13'd80,  13'd546,  
-13'd59,  -13'd28,  13'd703,  -13'd504,  -13'd408,  -13'd360,  13'd10,  -13'd42,  13'd93,  13'd381,  13'd143,  -13'd171,  -13'd128,  13'd115,  13'd270,  -13'd415,  
13'd560,  13'd368,  13'd231,  13'd161,  -13'd172,  -13'd390,  -13'd704,  -13'd976,  -13'd105,  -13'd21,  -13'd401,  -13'd160,  -13'd652,  13'd577,  13'd169,  13'd117,  
-13'd21,  -13'd197,  -13'd678,  -13'd67,  -13'd738,  13'd615,  13'd1,  -13'd92,  13'd560,  -13'd520,  13'd333,  -13'd99,  13'd173,  13'd149,  13'd330,  -13'd437,  
13'd550,  -13'd273,  13'd292,  13'd416,  13'd271,  -13'd149,  13'd146,  -13'd3,  13'd107,  -13'd455,  -13'd703,  13'd309,  13'd988,  13'd248,  13'd70,  13'd362,  
13'd181,  13'd704,  13'd21,  13'd11,  13'd650,  13'd7,  13'd148,  13'd329,  -13'd54,  13'd197,  13'd758,  13'd640,  -13'd60,  13'd844,  -13'd232,  -13'd216,  
-13'd21,  13'd268,  -13'd141,  -13'd84,  -13'd167,  13'd381,  13'd12,  13'd515,  -13'd888,  -13'd412,  -13'd55,  13'd295,  -13'd120,  13'd179,  -13'd70,  -13'd202,  
13'd1139,  13'd480,  13'd51,  13'd448,  -13'd84,  -13'd147,  13'd242,  13'd336,  -13'd498,  -13'd1133,  -13'd74,  -13'd51,  13'd33,  13'd336,  13'd469,  -13'd577,  
13'd174,  -13'd6,  -13'd907,  -13'd551,  -13'd375,  13'd199,  -13'd137,  -13'd193,  13'd518,  -13'd509,  -13'd304,  -13'd307,  13'd501,  13'd240,  -13'd49,  13'd747,  
13'd89,  13'd404,  -13'd42,  -13'd309,  13'd889,  13'd272,  -13'd135,  13'd251,  -13'd642,  -13'd143,  13'd136,  -13'd20,  -13'd10,  13'd629,  -13'd5,  13'd630,  
-13'd169,  -13'd370,  -13'd320,  -13'd188,  13'd1082,  -13'd849,  -13'd147,  13'd166,  -13'd180,  -13'd207,  -13'd87,  -13'd91,  13'd541,  -13'd382,  -13'd388,  -13'd28,  
13'd339,  13'd620,  -13'd663,  13'd8,  13'd54,  -13'd44,  13'd316,  -13'd203,  13'd497,  -13'd18,  -13'd847,  13'd86,  -13'd528,  13'd403,  -13'd586,  13'd596,  
13'd80,  -13'd150,  13'd103,  -13'd244,  -13'd320,  13'd229,  -13'd469,  13'd355,  -13'd378,  -13'd121,  -13'd587,  -13'd59,  13'd586,  13'd132,  -13'd526,  -13'd130,  
13'd1,  -13'd684,  -13'd340,  -13'd216,  -13'd484,  -13'd466,  13'd628,  -13'd589,  -13'd208,  -13'd854,  13'd257,  13'd469,  13'd562,  -13'd96,  13'd8,  13'd304,  
13'd220,  13'd640,  13'd716,  13'd107,  -13'd518,  13'd199,  -13'd726,  13'd407,  -13'd1230,  -13'd95,  13'd364,  -13'd11,  13'd294,  -13'd489,  -13'd167,  -13'd106,  
-13'd654,  -13'd425,  13'd32,  -13'd669,  13'd474,  -13'd616,  13'd481,  13'd386,  13'd550,  -13'd892,  -13'd709,  13'd52,  13'd331,  13'd425,  -13'd767,  -13'd194,  
-13'd1034,  -13'd180,  -13'd466,  -13'd408,  -13'd96,  13'd320,  -13'd174,  13'd420,  13'd330,  -13'd678,  -13'd289,  -13'd407,  -13'd206,  13'd920,  13'd157,  13'd175,  
-13'd639,  -13'd621,  13'd573,  -13'd112,  13'd188,  -13'd566,  13'd367,  -13'd164,  -13'd264,  -13'd201,  -13'd838,  -13'd375,  13'd88,  13'd733,  -13'd557,  13'd17,  
13'd22,  -13'd157,  -13'd749,  13'd41,  13'd198,  -13'd12,  13'd1,  13'd551,  -13'd933,  -13'd49,  -13'd478,  13'd148,  13'd346,  -13'd491,  13'd67,  -13'd238,  

13'd306,  13'd411,  13'd280,  13'd73,  -13'd403,  13'd68,  -13'd844,  -13'd4,  13'd376,  -13'd463,  -13'd613,  13'd551,  13'd436,  -13'd191,  -13'd403,  13'd380,  
13'd29,  -13'd91,  -13'd118,  13'd466,  -13'd92,  -13'd201,  -13'd609,  -13'd94,  -13'd101,  13'd368,  13'd523,  13'd149,  13'd506,  13'd1218,  -13'd721,  -13'd797,  
-13'd616,  13'd607,  13'd267,  -13'd393,  -13'd432,  13'd15,  -13'd636,  -13'd462,  13'd694,  -13'd249,  -13'd326,  -13'd130,  -13'd406,  13'd585,  13'd290,  -13'd79,  
13'd28,  13'd121,  -13'd124,  13'd204,  -13'd463,  13'd140,  -13'd590,  13'd124,  -13'd246,  -13'd262,  -13'd672,  13'd29,  -13'd468,  13'd383,  13'd853,  13'd378,  
13'd660,  13'd191,  -13'd785,  13'd853,  13'd354,  -13'd261,  -13'd198,  13'd219,  13'd556,  13'd346,  13'd262,  13'd94,  13'd578,  13'd611,  13'd565,  13'd251,  
13'd419,  -13'd631,  13'd272,  13'd406,  -13'd854,  13'd595,  -13'd391,  13'd681,  -13'd115,  13'd125,  -13'd743,  13'd80,  -13'd48,  13'd346,  13'd160,  13'd96,  
-13'd242,  -13'd1089,  13'd823,  -13'd227,  13'd229,  13'd311,  13'd484,  -13'd161,  -13'd259,  -13'd318,  13'd268,  -13'd453,  13'd7,  13'd481,  13'd704,  13'd222,  
13'd376,  -13'd39,  -13'd64,  -13'd94,  -13'd494,  13'd245,  13'd189,  -13'd620,  -13'd209,  13'd575,  -13'd545,  -13'd156,  -13'd617,  13'd940,  13'd329,  -13'd716,  
-13'd136,  13'd275,  -13'd87,  -13'd85,  13'd39,  -13'd365,  13'd42,  -13'd141,  13'd560,  -13'd203,  13'd141,  13'd564,  -13'd405,  -13'd694,  13'd2,  -13'd241,  
13'd420,  13'd563,  -13'd245,  -13'd217,  -13'd804,  13'd726,  -13'd251,  -13'd348,  13'd901,  13'd16,  13'd410,  13'd106,  13'd147,  13'd856,  -13'd534,  13'd948,  
-13'd30,  13'd122,  -13'd6,  13'd816,  -13'd478,  13'd307,  13'd19,  13'd407,  13'd153,  13'd476,  13'd733,  -13'd198,  13'd137,  -13'd339,  13'd131,  -13'd98,  
13'd165,  13'd612,  13'd1,  13'd299,  13'd343,  13'd243,  -13'd43,  13'd576,  -13'd221,  13'd576,  -13'd405,  -13'd263,  -13'd291,  13'd662,  -13'd47,  13'd499,  
-13'd603,  13'd32,  -13'd120,  -13'd801,  13'd644,  13'd304,  13'd368,  13'd13,  -13'd428,  -13'd135,  13'd353,  -13'd305,  -13'd302,  13'd220,  -13'd333,  13'd58,  
-13'd886,  13'd624,  -13'd174,  -13'd323,  13'd417,  -13'd513,  -13'd266,  -13'd115,  -13'd564,  -13'd57,  -13'd335,  13'd800,  -13'd907,  -13'd226,  13'd543,  13'd435,  
-13'd397,  13'd450,  13'd339,  13'd402,  13'd112,  13'd290,  13'd135,  13'd425,  13'd254,  -13'd76,  -13'd368,  -13'd249,  -13'd674,  -13'd22,  -13'd238,  -13'd79,  
-13'd237,  13'd543,  13'd521,  13'd54,  13'd38,  13'd369,  13'd361,  13'd672,  13'd150,  -13'd282,  -13'd11,  13'd324,  13'd480,  -13'd712,  13'd253,  -13'd64,  
13'd304,  13'd160,  13'd169,  -13'd404,  13'd760,  -13'd395,  -13'd178,  -13'd164,  -13'd266,  13'd412,  13'd26,  13'd138,  13'd144,  13'd65,  13'd699,  -13'd295,  
13'd216,  -13'd96,  -13'd410,  -13'd52,  13'd126,  13'd49,  -13'd474,  13'd246,  -13'd889,  -13'd495,  13'd839,  13'd135,  13'd397,  13'd587,  -13'd520,  -13'd142,  
13'd181,  13'd501,  13'd253,  13'd575,  13'd480,  13'd290,  13'd15,  13'd823,  13'd315,  -13'd241,  -13'd96,  13'd490,  13'd222,  13'd269,  -13'd49,  -13'd45,  
13'd1003,  13'd113,  -13'd203,  13'd376,  -13'd345,  -13'd52,  -13'd672,  13'd363,  13'd473,  13'd242,  -13'd2,  -13'd207,  -13'd392,  13'd406,  13'd149,  -13'd133,  
-13'd655,  13'd271,  -13'd617,  -13'd352,  -13'd700,  13'd456,  13'd1042,  13'd42,  13'd630,  -13'd376,  13'd17,  -13'd221,  -13'd570,  -13'd153,  -13'd32,  13'd549,  
-13'd512,  -13'd316,  -13'd187,  -13'd495,  13'd349,  13'd750,  13'd212,  13'd211,  13'd133,  13'd48,  13'd575,  13'd35,  13'd546,  -13'd662,  13'd842,  -13'd173,  
13'd485,  -13'd159,  -13'd953,  -13'd835,  13'd265,  -13'd39,  -13'd254,  13'd47,  13'd57,  13'd254,  13'd113,  13'd510,  13'd68,  13'd152,  -13'd629,  -13'd544,  
13'd1134,  13'd940,  13'd71,  13'd207,  13'd604,  13'd58,  13'd34,  13'd79,  -13'd202,  13'd749,  13'd309,  13'd356,  -13'd11,  13'd609,  13'd623,  -13'd88,  
-13'd447,  13'd785,  -13'd284,  13'd492,  -13'd274,  13'd199,  13'd481,  13'd978,  13'd437,  -13'd718,  -13'd406,  13'd884,  -13'd152,  -13'd476,  13'd313,  13'd557,  

-13'd272,  13'd472,  -13'd365,  -13'd136,  13'd569,  13'd377,  -13'd133,  13'd220,  13'd244,  -13'd18,  -13'd721,  -13'd137,  13'd174,  13'd282,  -13'd598,  13'd631,  
13'd412,  13'd401,  -13'd617,  -13'd350,  13'd114,  13'd283,  13'd48,  13'd352,  -13'd805,  -13'd362,  -13'd417,  -13'd445,  13'd158,  13'd103,  -13'd408,  -13'd472,  
-13'd494,  13'd431,  -13'd126,  13'd580,  -13'd387,  -13'd58,  13'd238,  -13'd45,  13'd167,  -13'd28,  -13'd25,  -13'd184,  13'd66,  13'd624,  13'd461,  -13'd624,  
13'd524,  -13'd44,  -13'd552,  -13'd339,  -13'd228,  13'd116,  13'd384,  -13'd528,  13'd39,  13'd341,  13'd310,  -13'd725,  -13'd352,  13'd158,  13'd28,  -13'd39,  
13'd305,  -13'd374,  13'd692,  13'd172,  13'd376,  -13'd523,  -13'd199,  13'd107,  -13'd602,  13'd132,  -13'd512,  -13'd261,  -13'd39,  -13'd625,  -13'd147,  13'd478,  
13'd65,  -13'd229,  13'd505,  -13'd12,  -13'd289,  -13'd141,  13'd327,  -13'd398,  -13'd29,  -13'd253,  13'd35,  13'd103,  -13'd306,  -13'd226,  13'd260,  -13'd78,  
-13'd174,  -13'd26,  -13'd476,  13'd301,  13'd138,  -13'd23,  -13'd165,  -13'd172,  -13'd345,  13'd230,  13'd186,  13'd449,  -13'd545,  13'd654,  -13'd121,  -13'd312,  
13'd62,  -13'd193,  13'd47,  -13'd880,  13'd275,  -13'd14,  13'd78,  -13'd771,  13'd191,  -13'd14,  -13'd310,  13'd140,  -13'd572,  13'd240,  13'd142,  -13'd352,  
-13'd43,  -13'd45,  13'd257,  13'd88,  13'd81,  -13'd693,  -13'd283,  -13'd335,  -13'd14,  -13'd336,  13'd154,  13'd127,  -13'd15,  13'd238,  13'd85,  13'd54,  
13'd185,  -13'd415,  13'd263,  13'd306,  13'd217,  13'd179,  -13'd292,  13'd149,  13'd710,  13'd175,  13'd121,  13'd32,  -13'd51,  13'd424,  -13'd263,  -13'd534,  
-13'd104,  -13'd434,  -13'd311,  13'd75,  -13'd236,  13'd257,  13'd331,  -13'd849,  -13'd90,  13'd264,  -13'd142,  13'd6,  13'd280,  13'd346,  13'd540,  -13'd584,  
13'd13,  -13'd43,  -13'd645,  -13'd168,  -13'd429,  -13'd521,  13'd490,  -13'd438,  -13'd780,  -13'd95,  13'd129,  -13'd221,  -13'd313,  13'd28,  -13'd721,  -13'd246,  
-13'd170,  13'd472,  13'd450,  13'd24,  -13'd312,  -13'd149,  -13'd395,  13'd212,  -13'd547,  -13'd793,  -13'd100,  13'd249,  13'd161,  13'd153,  -13'd615,  13'd398,  
-13'd154,  -13'd697,  13'd11,  -13'd236,  13'd89,  -13'd30,  13'd523,  -13'd534,  -13'd392,  -13'd246,  -13'd708,  13'd98,  -13'd324,  13'd539,  -13'd575,  -13'd504,  
-13'd302,  -13'd740,  -13'd269,  13'd1,  -13'd387,  13'd348,  -13'd327,  13'd167,  -13'd105,  -13'd530,  13'd132,  -13'd680,  -13'd458,  -13'd253,  13'd563,  13'd92,  
-13'd44,  13'd300,  13'd601,  -13'd565,  -13'd200,  13'd571,  -13'd771,  -13'd53,  -13'd641,  -13'd557,  13'd343,  -13'd635,  13'd145,  13'd649,  13'd343,  -13'd107,  
-13'd539,  -13'd447,  13'd118,  -13'd466,  -13'd517,  13'd15,  13'd683,  -13'd233,  13'd248,  13'd278,  13'd143,  13'd124,  -13'd101,  13'd580,  -13'd167,  13'd76,  
-13'd163,  13'd239,  -13'd517,  -13'd538,  13'd94,  -13'd60,  -13'd557,  13'd103,  -13'd170,  -13'd13,  13'd333,  13'd421,  -13'd450,  -13'd408,  -13'd517,  -13'd215,  
-13'd733,  -13'd190,  -13'd423,  13'd229,  13'd104,  13'd481,  -13'd62,  -13'd50,  -13'd176,  13'd182,  13'd297,  -13'd135,  -13'd109,  13'd88,  -13'd97,  -13'd398,  
-13'd414,  -13'd563,  13'd241,  13'd53,  13'd400,  13'd133,  13'd77,  -13'd97,  13'd201,  -13'd252,  -13'd693,  13'd313,  -13'd248,  13'd42,  -13'd368,  13'd207,  
-13'd55,  -13'd167,  13'd258,  13'd720,  13'd235,  -13'd403,  13'd227,  13'd10,  -13'd54,  13'd425,  13'd59,  -13'd13,  13'd99,  -13'd441,  -13'd433,  -13'd241,  
-13'd475,  -13'd69,  13'd634,  -13'd113,  -13'd176,  -13'd22,  -13'd496,  13'd32,  -13'd410,  13'd104,  13'd505,  -13'd84,  13'd106,  -13'd32,  -13'd161,  13'd327,  
-13'd187,  -13'd111,  13'd38,  -13'd168,  13'd233,  13'd381,  -13'd486,  13'd60,  13'd314,  -13'd442,  -13'd374,  -13'd642,  -13'd249,  -13'd749,  -13'd693,  -13'd99,  
-13'd164,  13'd679,  -13'd385,  13'd64,  -13'd175,  -13'd251,  13'd6,  13'd43,  13'd311,  13'd368,  -13'd455,  -13'd273,  -13'd849,  -13'd159,  -13'd380,  -13'd807,  
-13'd610,  13'd157,  -13'd235,  -13'd212,  -13'd680,  13'd285,  -13'd564,  13'd429,  -13'd316,  13'd535,  -13'd245,  -13'd462,  13'd13,  -13'd186,  -13'd768,  13'd106,  

-13'd280,  -13'd124,  13'd571,  -13'd537,  -13'd470,  13'd451,  13'd2,  -13'd567,  -13'd299,  13'd129,  13'd226,  -13'd203,  13'd75,  13'd556,  -13'd533,  -13'd384,  
-13'd93,  13'd91,  13'd443,  13'd256,  -13'd208,  -13'd34,  13'd343,  13'd267,  13'd285,  -13'd397,  -13'd37,  13'd635,  13'd254,  13'd538,  -13'd192,  -13'd89,  
13'd536,  13'd164,  13'd316,  13'd221,  13'd48,  13'd117,  13'd306,  -13'd39,  13'd137,  -13'd389,  -13'd132,  -13'd373,  13'd607,  -13'd128,  -13'd324,  13'd123,  
13'd728,  -13'd80,  -13'd633,  -13'd37,  -13'd467,  13'd147,  13'd631,  13'd269,  -13'd121,  -13'd645,  13'd76,  -13'd140,  13'd395,  -13'd1233,  -13'd420,  13'd623,  
13'd516,  13'd853,  -13'd374,  13'd574,  13'd47,  -13'd155,  13'd611,  -13'd211,  13'd230,  13'd173,  -13'd24,  13'd534,  13'd567,  13'd676,  13'd114,  13'd1228,  
13'd193,  13'd157,  13'd390,  -13'd58,  -13'd359,  13'd474,  -13'd144,  -13'd327,  -13'd162,  13'd174,  -13'd269,  13'd710,  13'd346,  13'd185,  -13'd324,  13'd706,  
-13'd323,  13'd346,  13'd313,  13'd573,  -13'd665,  13'd332,  13'd152,  13'd297,  13'd491,  -13'd723,  -13'd130,  13'd100,  -13'd414,  -13'd452,  -13'd253,  -13'd142,  
-13'd401,  13'd248,  -13'd364,  13'd75,  13'd696,  -13'd5,  -13'd260,  13'd668,  -13'd12,  13'd158,  -13'd475,  -13'd65,  13'd767,  -13'd264,  -13'd752,  -13'd170,  
13'd134,  13'd185,  -13'd806,  13'd345,  13'd335,  -13'd231,  -13'd744,  13'd198,  13'd167,  13'd759,  13'd740,  -13'd153,  13'd287,  -13'd1098,  13'd735,  13'd486,  
-13'd101,  -13'd1074,  -13'd393,  13'd924,  13'd803,  13'd473,  -13'd237,  -13'd217,  13'd45,  -13'd298,  13'd387,  13'd85,  13'd463,  13'd326,  13'd310,  13'd515,  
-13'd429,  13'd153,  -13'd164,  -13'd261,  -13'd890,  -13'd722,  13'd650,  13'd243,  13'd172,  13'd116,  -13'd996,  13'd96,  -13'd366,  13'd119,  13'd940,  13'd417,  
-13'd659,  13'd219,  -13'd211,  -13'd286,  -13'd106,  -13'd61,  13'd231,  13'd484,  13'd17,  13'd128,  -13'd361,  -13'd93,  -13'd896,  -13'd85,  13'd440,  -13'd563,  
-13'd455,  -13'd130,  13'd840,  13'd833,  -13'd502,  -13'd361,  13'd7,  -13'd35,  13'd360,  13'd725,  -13'd626,  -13'd361,  -13'd323,  13'd212,  13'd526,  -13'd132,  
-13'd225,  13'd179,  -13'd1048,  -13'd215,  13'd531,  13'd153,  13'd447,  13'd135,  -13'd380,  13'd49,  -13'd193,  -13'd334,  13'd863,  -13'd635,  13'd466,  13'd662,  
-13'd1236,  -13'd497,  13'd7,  -13'd164,  13'd517,  -13'd646,  -13'd598,  -13'd59,  13'd539,  13'd149,  13'd347,  -13'd386,  -13'd880,  -13'd304,  -13'd37,  13'd577,  
-13'd455,  13'd544,  13'd161,  13'd686,  -13'd184,  -13'd295,  -13'd248,  -13'd90,  -13'd330,  13'd69,  -13'd1367,  -13'd83,  13'd104,  -13'd51,  13'd319,  13'd129,  
-13'd286,  -13'd502,  13'd354,  13'd17,  13'd335,  13'd563,  13'd27,  -13'd174,  -13'd1148,  13'd330,  -13'd776,  -13'd417,  13'd756,  13'd20,  13'd227,  -13'd299,  
-13'd524,  13'd332,  13'd367,  -13'd239,  13'd526,  -13'd77,  -13'd384,  -13'd284,  -13'd516,  13'd293,  13'd681,  13'd753,  13'd178,  13'd960,  -13'd674,  13'd257,  
-13'd331,  -13'd379,  13'd460,  13'd291,  13'd225,  -13'd83,  13'd365,  -13'd483,  -13'd155,  -13'd105,  13'd1038,  -13'd359,  -13'd127,  -13'd427,  13'd117,  13'd229,  
13'd76,  13'd641,  13'd55,  -13'd192,  13'd463,  13'd273,  13'd280,  13'd16,  13'd338,  -13'd292,  -13'd308,  13'd265,  -13'd20,  13'd233,  13'd81,  13'd71,  
-13'd292,  13'd410,  -13'd906,  -13'd37,  -13'd338,  -13'd158,  13'd270,  13'd148,  13'd625,  13'd211,  -13'd671,  -13'd106,  -13'd161,  13'd25,  -13'd337,  -13'd545,  
13'd293,  13'd358,  13'd310,  -13'd184,  -13'd46,  -13'd301,  13'd284,  13'd203,  13'd31,  -13'd569,  -13'd397,  13'd924,  -13'd337,  -13'd151,  13'd296,  13'd139,  
-13'd705,  13'd477,  -13'd660,  -13'd236,  -13'd613,  -13'd491,  13'd740,  -13'd39,  13'd142,  13'd372,  -13'd223,  -13'd225,  13'd290,  13'd234,  13'd252,  -13'd9,  
13'd203,  -13'd19,  13'd33,  -13'd277,  -13'd349,  -13'd564,  13'd90,  13'd458,  13'd323,  -13'd511,  13'd481,  13'd198,  -13'd603,  13'd608,  -13'd99,  -13'd206,  
13'd698,  -13'd298,  -13'd807,  -13'd246,  13'd18,  13'd157,  13'd734,  13'd375,  -13'd318,  -13'd762,  -13'd8,  -13'd405,  -13'd412,  13'd982,  -13'd73,  -13'd742,  

-13'd638,  -13'd482,  -13'd834,  -13'd272,  -13'd221,  -13'd343,  13'd1360,  -13'd659,  13'd77,  13'd471,  -13'd191,  -13'd472,  -13'd284,  -13'd418,  -13'd621,  -13'd549,  
13'd156,  -13'd558,  13'd82,  13'd77,  -13'd237,  13'd6,  13'd118,  13'd122,  13'd732,  13'd336,  -13'd129,  -13'd340,  -13'd237,  13'd401,  -13'd874,  13'd30,  
13'd440,  13'd139,  -13'd441,  -13'd826,  13'd183,  -13'd76,  -13'd476,  -13'd402,  13'd175,  -13'd434,  13'd226,  -13'd656,  13'd366,  -13'd227,  -13'd17,  13'd375,  
13'd466,  13'd546,  13'd232,  13'd322,  13'd444,  13'd210,  -13'd481,  -13'd53,  13'd205,  13'd620,  13'd68,  13'd121,  -13'd263,  -13'd206,  13'd698,  -13'd26,  
-13'd1014,  -13'd173,  13'd770,  13'd195,  13'd116,  13'd53,  -13'd94,  -13'd33,  -13'd556,  13'd763,  -13'd4,  -13'd36,  -13'd61,  -13'd261,  13'd290,  -13'd353,  
-13'd407,  13'd49,  13'd671,  13'd179,  -13'd533,  13'd211,  13'd144,  -13'd243,  -13'd235,  -13'd361,  13'd102,  -13'd110,  -13'd593,  -13'd449,  -13'd30,  -13'd113,  
13'd439,  13'd281,  -13'd293,  13'd879,  -13'd728,  13'd730,  -13'd644,  -13'd862,  13'd440,  -13'd85,  13'd216,  -13'd232,  13'd15,  -13'd721,  -13'd761,  -13'd198,  
-13'd18,  -13'd182,  13'd84,  13'd176,  13'd274,  -13'd280,  13'd144,  -13'd577,  -13'd101,  -13'd296,  13'd702,  -13'd207,  13'd437,  -13'd360,  -13'd478,  13'd813,  
-13'd577,  13'd519,  13'd194,  13'd320,  13'd283,  -13'd335,  13'd99,  13'd188,  -13'd158,  13'd207,  13'd86,  -13'd597,  -13'd230,  13'd420,  -13'd306,  13'd196,  
-13'd51,  -13'd159,  13'd803,  13'd257,  13'd217,  13'd591,  -13'd279,  13'd273,  -13'd192,  13'd323,  -13'd708,  13'd620,  -13'd415,  13'd202,  -13'd90,  -13'd781,  
13'd394,  13'd571,  -13'd384,  13'd597,  -13'd1484,  -13'd672,  13'd338,  13'd47,  13'd7,  13'd103,  -13'd818,  13'd234,  13'd38,  -13'd411,  -13'd113,  -13'd18,  
13'd254,  13'd160,  13'd291,  -13'd129,  -13'd510,  -13'd213,  13'd341,  13'd259,  13'd1237,  -13'd430,  13'd459,  -13'd457,  13'd93,  13'd572,  -13'd197,  13'd330,  
-13'd545,  13'd397,  -13'd81,  13'd394,  13'd913,  -13'd290,  13'd504,  13'd121,  13'd266,  13'd49,  13'd13,  13'd138,  13'd83,  -13'd53,  -13'd594,  -13'd307,  
13'd672,  -13'd213,  -13'd257,  -13'd159,  13'd261,  -13'd521,  -13'd201,  13'd522,  -13'd891,  -13'd90,  13'd257,  13'd368,  -13'd394,  13'd394,  13'd653,  -13'd584,  
13'd102,  13'd141,  13'd654,  13'd234,  13'd155,  13'd156,  -13'd182,  13'd323,  13'd780,  13'd183,  13'd138,  13'd102,  13'd656,  13'd386,  13'd578,  13'd230,  
-13'd34,  -13'd271,  13'd387,  13'd18,  -13'd479,  -13'd63,  13'd383,  13'd258,  13'd100,  -13'd183,  -13'd143,  13'd337,  13'd113,  13'd619,  13'd644,  -13'd478,  
13'd108,  13'd231,  13'd211,  13'd488,  -13'd405,  13'd120,  13'd198,  13'd39,  13'd544,  -13'd442,  13'd526,  -13'd95,  -13'd471,  -13'd260,  -13'd326,  -13'd543,  
-13'd521,  -13'd649,  -13'd565,  -13'd355,  -13'd20,  13'd675,  13'd417,  -13'd660,  -13'd105,  13'd361,  13'd897,  -13'd280,  -13'd245,  -13'd485,  -13'd160,  13'd413,  
-13'd486,  13'd590,  -13'd383,  -13'd471,  13'd41,  13'd563,  13'd128,  -13'd94,  -13'd253,  13'd677,  13'd135,  -13'd214,  13'd766,  13'd132,  -13'd151,  13'd11,  
13'd133,  -13'd191,  13'd176,  13'd39,  13'd476,  13'd641,  -13'd617,  13'd403,  13'd158,  13'd406,  13'd68,  13'd282,  13'd423,  -13'd601,  13'd587,  13'd1110,  
-13'd225,  -13'd676,  13'd599,  13'd187,  13'd509,  -13'd170,  -13'd866,  13'd584,  -13'd14,  -13'd316,  13'd20,  -13'd12,  -13'd216,  13'd804,  13'd753,  -13'd96,  
-13'd963,  -13'd450,  -13'd115,  13'd288,  13'd16,  13'd355,  -13'd100,  13'd587,  -13'd304,  -13'd365,  13'd204,  -13'd52,  13'd259,  -13'd398,  13'd9,  -13'd509,  
-13'd376,  -13'd1425,  -13'd301,  13'd238,  13'd136,  13'd384,  -13'd561,  -13'd419,  -13'd638,  -13'd78,  13'd376,  -13'd404,  13'd75,  -13'd614,  -13'd130,  13'd626,  
-13'd215,  13'd128,  13'd122,  -13'd618,  13'd451,  -13'd518,  13'd125,  13'd95,  13'd75,  13'd897,  13'd290,  13'd174,  -13'd252,  -13'd615,  13'd253,  -13'd338,  
-13'd761,  13'd133,  -13'd629,  -13'd648,  13'd508,  -13'd732,  -13'd462,  -13'd217,  13'd648,  13'd1130,  -13'd171,  13'd195,  13'd458,  -13'd1055,  13'd8,  -13'd358,  

-13'd619,  -13'd482,  13'd138,  -13'd318,  -13'd715,  13'd143,  -13'd877,  -13'd225,  -13'd538,  -13'd265,  -13'd391,  -13'd483,  13'd223,  13'd708,  13'd322,  13'd113,  
13'd7,  -13'd63,  13'd4,  -13'd454,  13'd0,  13'd107,  -13'd99,  13'd435,  -13'd539,  13'd872,  -13'd185,  -13'd289,  13'd618,  -13'd199,  -13'd712,  13'd360,  
-13'd322,  -13'd624,  13'd19,  -13'd444,  13'd75,  13'd504,  -13'd90,  13'd576,  13'd240,  -13'd192,  -13'd246,  -13'd16,  13'd781,  -13'd300,  13'd418,  -13'd306,  
-13'd254,  13'd875,  13'd79,  13'd225,  13'd71,  -13'd142,  -13'd794,  -13'd162,  -13'd204,  -13'd485,  13'd418,  -13'd70,  -13'd119,  -13'd1036,  13'd835,  -13'd746,  
13'd858,  -13'd38,  -13'd32,  13'd998,  -13'd78,  -13'd89,  -13'd11,  -13'd180,  -13'd368,  -13'd122,  13'd500,  13'd370,  -13'd404,  -13'd255,  13'd586,  -13'd372,  
-13'd542,  -13'd336,  13'd68,  -13'd898,  -13'd328,  13'd327,  13'd138,  -13'd608,  13'd256,  -13'd378,  -13'd510,  -13'd134,  13'd23,  -13'd293,  13'd404,  13'd636,  
13'd756,  -13'd272,  13'd108,  13'd439,  -13'd277,  -13'd313,  13'd53,  13'd31,  -13'd485,  -13'd68,  -13'd2,  -13'd216,  13'd339,  13'd129,  13'd19,  13'd104,  
13'd1113,  13'd320,  13'd107,  13'd66,  13'd9,  13'd329,  13'd1407,  13'd32,  13'd138,  -13'd450,  -13'd872,  -13'd425,  -13'd182,  -13'd40,  13'd383,  -13'd994,  
13'd586,  13'd693,  13'd449,  13'd303,  13'd786,  13'd9,  -13'd71,  -13'd341,  13'd944,  13'd487,  13'd446,  13'd767,  -13'd156,  13'd731,  13'd748,  -13'd92,  
13'd85,  -13'd470,  -13'd80,  -13'd168,  -13'd393,  13'd271,  13'd342,  13'd427,  13'd881,  -13'd63,  13'd384,  13'd843,  -13'd240,  13'd294,  13'd44,  -13'd528,  
-13'd859,  -13'd149,  -13'd193,  13'd96,  -13'd1013,  13'd217,  13'd202,  -13'd385,  -13'd551,  -13'd763,  -13'd310,  13'd100,  -13'd405,  13'd864,  13'd437,  -13'd96,  
13'd1097,  13'd228,  -13'd71,  -13'd377,  -13'd532,  -13'd92,  -13'd35,  -13'd374,  -13'd100,  -13'd203,  -13'd47,  13'd777,  13'd125,  13'd162,  -13'd612,  13'd305,  
13'd385,  13'd814,  13'd375,  -13'd308,  13'd499,  13'd24,  13'd923,  -13'd45,  13'd217,  13'd98,  -13'd258,  13'd331,  13'd141,  13'd374,  13'd130,  -13'd142,  
13'd446,  13'd470,  13'd276,  -13'd248,  -13'd254,  13'd377,  -13'd150,  13'd27,  -13'd153,  -13'd811,  13'd752,  13'd355,  -13'd350,  -13'd102,  13'd519,  13'd352,  
13'd228,  13'd442,  -13'd150,  -13'd211,  -13'd304,  -13'd56,  -13'd96,  -13'd0,  13'd1022,  -13'd291,  13'd451,  -13'd335,  -13'd88,  13'd731,  -13'd29,  -13'd630,  
13'd90,  -13'd243,  -13'd48,  13'd107,  -13'd294,  -13'd352,  13'd584,  -13'd516,  -13'd628,  -13'd282,  -13'd56,  13'd574,  13'd242,  -13'd52,  13'd230,  -13'd35,  
13'd851,  13'd535,  13'd254,  -13'd167,  -13'd305,  -13'd509,  13'd340,  13'd85,  -13'd684,  -13'd650,  -13'd266,  -13'd42,  13'd430,  -13'd137,  -13'd580,  13'd95,  
13'd418,  13'd220,  -13'd491,  13'd41,  -13'd660,  -13'd346,  13'd466,  -13'd220,  -13'd706,  -13'd385,  13'd778,  -13'd192,  -13'd160,  13'd705,  -13'd699,  -13'd470,  
13'd294,  13'd308,  13'd678,  -13'd96,  -13'd629,  13'd329,  13'd485,  13'd150,  -13'd228,  -13'd761,  13'd684,  -13'd1,  13'd151,  -13'd545,  13'd47,  13'd274,  
-13'd458,  -13'd368,  -13'd869,  -13'd973,  -13'd176,  -13'd851,  13'd322,  13'd157,  -13'd814,  -13'd1604,  -13'd111,  -13'd905,  13'd296,  13'd180,  -13'd1089,  -13'd76,  
-13'd337,  13'd191,  -13'd136,  -13'd138,  -13'd815,  -13'd36,  -13'd171,  13'd446,  -13'd488,  13'd323,  13'd536,  13'd381,  -13'd4,  13'd538,  13'd420,  -13'd64,  
13'd510,  -13'd246,  13'd836,  13'd159,  -13'd215,  -13'd152,  13'd353,  -13'd3,  -13'd584,  13'd274,  -13'd68,  -13'd495,  13'd218,  13'd316,  13'd192,  13'd352,  
-13'd552,  13'd563,  13'd116,  -13'd582,  13'd156,  -13'd1130,  13'd645,  -13'd151,  -13'd366,  13'd1039,  -13'd311,  -13'd686,  -13'd103,  13'd780,  -13'd507,  -13'd460,  
-13'd981,  -13'd974,  13'd62,  -13'd1619,  -13'd416,  -13'd737,  13'd68,  -13'd54,  13'd13,  -13'd430,  -13'd644,  -13'd1049,  -13'd546,  -13'd26,  -13'd685,  -13'd389,  
13'd107,  -13'd671,  -13'd846,  -13'd1158,  -13'd1082,  -13'd780,  -13'd614,  -13'd380,  -13'd651,  -13'd1258,  -13'd423,  -13'd1208,  -13'd1444,  -13'd373,  -13'd707,  -13'd1244,  

-13'd114,  13'd280,  13'd461,  13'd183,  -13'd382,  -13'd298,  -13'd68,  -13'd222,  13'd336,  -13'd125,  13'd130,  -13'd194,  13'd376,  13'd200,  -13'd277,  13'd582,  
13'd149,  13'd851,  13'd1282,  13'd228,  13'd210,  -13'd322,  13'd490,  13'd172,  13'd562,  -13'd208,  13'd502,  13'd271,  13'd155,  13'd32,  -13'd337,  -13'd179,  
-13'd258,  13'd90,  13'd698,  -13'd117,  13'd461,  13'd757,  13'd776,  13'd277,  -13'd117,  -13'd1186,  -13'd169,  13'd541,  -13'd263,  13'd1553,  13'd428,  -13'd25,  
13'd535,  13'd17,  13'd63,  13'd204,  13'd481,  -13'd371,  -13'd323,  13'd494,  13'd248,  13'd747,  13'd337,  13'd399,  -13'd560,  13'd591,  13'd92,  13'd553,  
-13'd816,  -13'd367,  -13'd3,  13'd546,  -13'd1301,  -13'd212,  -13'd366,  13'd393,  13'd65,  13'd518,  -13'd472,  13'd381,  -13'd649,  -13'd541,  13'd94,  -13'd501,  
-13'd336,  13'd888,  13'd508,  13'd195,  13'd406,  -13'd310,  13'd496,  -13'd71,  -13'd818,  -13'd536,  13'd74,  -13'd615,  -13'd493,  13'd584,  -13'd236,  -13'd298,  
13'd330,  -13'd199,  13'd153,  -13'd562,  13'd9,  13'd34,  13'd360,  -13'd568,  13'd17,  13'd257,  13'd1121,  13'd39,  13'd546,  13'd893,  13'd172,  13'd111,  
-13'd338,  -13'd89,  13'd147,  13'd175,  -13'd446,  13'd381,  13'd168,  -13'd839,  13'd25,  -13'd227,  13'd216,  13'd15,  13'd471,  13'd247,  -13'd250,  13'd608,  
-13'd257,  13'd1003,  -13'd539,  13'd272,  13'd1002,  13'd44,  -13'd689,  -13'd124,  -13'd193,  13'd203,  -13'd1,  13'd255,  -13'd521,  -13'd488,  13'd159,  -13'd671,  
13'd445,  -13'd994,  13'd206,  -13'd27,  13'd280,  -13'd160,  13'd10,  -13'd529,  -13'd73,  13'd708,  -13'd77,  13'd14,  -13'd540,  13'd199,  13'd287,  -13'd335,  
13'd291,  13'd360,  13'd151,  -13'd878,  -13'd983,  -13'd973,  13'd1081,  -13'd643,  -13'd907,  -13'd596,  13'd738,  13'd365,  -13'd1036,  13'd625,  13'd299,  13'd261,  
13'd362,  -13'd187,  13'd690,  -13'd563,  -13'd456,  13'd126,  13'd532,  -13'd112,  13'd41,  -13'd150,  -13'd198,  -13'd216,  -13'd742,  13'd43,  -13'd308,  -13'd294,  
-13'd184,  13'd676,  -13'd397,  -13'd1109,  13'd488,  -13'd628,  13'd176,  13'd290,  13'd662,  -13'd55,  -13'd358,  -13'd187,  -13'd495,  13'd151,  13'd381,  -13'd41,  
-13'd367,  13'd865,  -13'd175,  13'd341,  -13'd96,  -13'd454,  13'd575,  13'd282,  -13'd310,  -13'd487,  13'd134,  -13'd237,  -13'd358,  13'd173,  13'd192,  -13'd308,  
-13'd813,  13'd156,  13'd114,  -13'd474,  -13'd411,  -13'd454,  13'd235,  -13'd204,  13'd58,  -13'd722,  -13'd626,  -13'd15,  -13'd677,  -13'd370,  13'd363,  13'd307,  
13'd2,  -13'd348,  13'd499,  -13'd355,  -13'd392,  13'd454,  13'd224,  13'd331,  -13'd421,  13'd197,  13'd5,  -13'd214,  -13'd348,  13'd703,  -13'd319,  -13'd248,  
13'd370,  -13'd124,  13'd255,  -13'd1026,  -13'd396,  -13'd0,  -13'd324,  -13'd256,  13'd291,  -13'd179,  -13'd268,  13'd33,  -13'd958,  13'd153,  -13'd371,  -13'd565,  
13'd695,  -13'd388,  13'd524,  13'd508,  -13'd387,  13'd276,  13'd155,  13'd751,  -13'd890,  -13'd128,  13'd395,  13'd486,  13'd208,  13'd834,  13'd665,  -13'd446,  
-13'd494,  13'd111,  -13'd597,  13'd1001,  -13'd589,  -13'd1,  -13'd538,  -13'd22,  13'd82,  13'd122,  -13'd708,  -13'd407,  13'd17,  -13'd277,  13'd350,  -13'd490,  
13'd729,  -13'd27,  13'd642,  -13'd64,  13'd42,  13'd156,  13'd276,  -13'd269,  13'd374,  13'd482,  13'd16,  13'd735,  13'd251,  -13'd515,  -13'd174,  13'd337,  
13'd23,  -13'd777,  13'd861,  -13'd501,  -13'd780,  -13'd662,  -13'd713,  -13'd303,  -13'd592,  13'd819,  -13'd1240,  13'd939,  -13'd68,  13'd671,  13'd325,  -13'd399,  
13'd94,  13'd656,  13'd785,  -13'd460,  -13'd293,  13'd16,  -13'd572,  13'd797,  13'd543,  13'd385,  -13'd693,  13'd377,  13'd123,  13'd140,  13'd202,  13'd145,  
13'd267,  13'd345,  13'd23,  13'd916,  13'd296,  13'd1187,  -13'd362,  13'd1031,  13'd540,  -13'd966,  -13'd350,  -13'd1031,  13'd560,  -13'd516,  13'd49,  13'd168,  
-13'd439,  -13'd481,  13'd356,  -13'd456,  13'd362,  -13'd290,  -13'd591,  -13'd78,  -13'd757,  13'd379,  13'd655,  -13'd977,  -13'd156,  -13'd509,  13'd243,  13'd299,  
-13'd139,  -13'd831,  -13'd558,  13'd604,  13'd930,  -13'd544,  -13'd334,  13'd673,  13'd161,  13'd1256,  13'd720,  13'd414,  -13'd219,  13'd28,  13'd235,  13'd881,  

13'd177,  13'd292,  13'd164,  13'd236,  13'd33,  13'd83,  -13'd759,  13'd36,  13'd98,  -13'd634,  13'd299,  -13'd87,  -13'd13,  -13'd447,  -13'd43,  13'd275,  
13'd526,  -13'd42,  -13'd271,  -13'd493,  13'd382,  13'd702,  13'd37,  -13'd103,  -13'd291,  -13'd242,  -13'd547,  13'd313,  13'd672,  -13'd239,  13'd337,  13'd313,  
13'd199,  -13'd164,  13'd57,  13'd335,  13'd95,  13'd437,  -13'd82,  -13'd488,  13'd320,  13'd531,  -13'd789,  -13'd584,  -13'd438,  13'd390,  13'd248,  13'd266,  
-13'd582,  -13'd137,  -13'd579,  -13'd180,  -13'd283,  -13'd120,  -13'd196,  -13'd100,  13'd772,  13'd465,  -13'd114,  -13'd40,  -13'd33,  13'd1009,  13'd670,  -13'd3,  
-13'd698,  -13'd344,  -13'd248,  13'd167,  13'd197,  -13'd12,  -13'd688,  13'd287,  13'd568,  13'd438,  13'd348,  13'd156,  -13'd590,  13'd189,  13'd357,  -13'd223,  
13'd187,  13'd54,  -13'd1026,  13'd208,  -13'd323,  -13'd315,  -13'd340,  -13'd776,  13'd414,  13'd810,  13'd304,  13'd111,  13'd436,  -13'd735,  -13'd351,  -13'd128,  
-13'd37,  -13'd4,  -13'd173,  -13'd533,  13'd420,  13'd140,  -13'd660,  -13'd174,  -13'd693,  13'd487,  -13'd195,  -13'd242,  -13'd21,  13'd237,  13'd86,  13'd297,  
-13'd604,  13'd1135,  13'd286,  -13'd144,  13'd36,  -13'd251,  13'd231,  -13'd431,  13'd590,  13'd739,  -13'd201,  13'd868,  -13'd356,  13'd688,  -13'd423,  13'd567,  
13'd64,  -13'd522,  13'd431,  13'd288,  -13'd130,  13'd65,  -13'd529,  -13'd146,  -13'd420,  -13'd813,  -13'd742,  13'd317,  -13'd17,  13'd551,  13'd229,  13'd484,  
-13'd291,  13'd429,  13'd664,  -13'd670,  -13'd62,  13'd441,  13'd463,  -13'd305,  13'd79,  13'd145,  13'd159,  13'd564,  -13'd124,  13'd230,  -13'd320,  -13'd307,  
-13'd485,  13'd8,  13'd198,  -13'd234,  -13'd579,  -13'd4,  13'd70,  -13'd883,  13'd266,  -13'd309,  13'd353,  13'd8,  -13'd1029,  -13'd828,  -13'd681,  13'd415,  
13'd622,  13'd478,  -13'd333,  13'd105,  -13'd244,  13'd805,  13'd501,  -13'd54,  13'd957,  -13'd81,  -13'd697,  13'd10,  -13'd219,  13'd213,  -13'd642,  -13'd361,  
13'd273,  13'd575,  -13'd528,  -13'd247,  13'd557,  -13'd73,  -13'd430,  13'd201,  13'd22,  -13'd217,  -13'd688,  13'd845,  13'd698,  -13'd129,  13'd60,  -13'd602,  
-13'd254,  13'd27,  13'd372,  13'd335,  -13'd118,  -13'd472,  13'd474,  -13'd659,  13'd246,  13'd165,  -13'd49,  -13'd62,  13'd2,  13'd230,  -13'd135,  13'd222,  
13'd339,  13'd46,  -13'd707,  13'd357,  13'd638,  13'd165,  -13'd231,  -13'd501,  -13'd391,  13'd59,  -13'd694,  13'd547,  13'd374,  -13'd753,  -13'd386,  -13'd129,  
13'd418,  -13'd709,  13'd456,  13'd432,  -13'd305,  -13'd53,  13'd718,  13'd57,  13'd482,  13'd14,  13'd511,  13'd81,  -13'd331,  13'd301,  13'd22,  13'd66,  
13'd129,  -13'd497,  -13'd123,  13'd382,  13'd157,  13'd723,  13'd554,  13'd400,  13'd86,  13'd110,  13'd338,  13'd425,  -13'd230,  13'd286,  13'd419,  13'd32,  
13'd521,  13'd43,  -13'd459,  13'd700,  -13'd94,  13'd133,  13'd111,  -13'd61,  -13'd751,  13'd533,  13'd52,  13'd20,  13'd371,  -13'd558,  13'd519,  -13'd299,  
-13'd158,  -13'd709,  -13'd548,  13'd155,  13'd428,  13'd131,  13'd157,  13'd227,  -13'd48,  -13'd242,  13'd511,  13'd483,  -13'd343,  -13'd663,  13'd788,  -13'd293,  
-13'd109,  13'd38,  -13'd547,  13'd124,  13'd199,  13'd479,  -13'd142,  13'd21,  -13'd342,  13'd524,  13'd741,  13'd423,  -13'd197,  -13'd330,  13'd729,  13'd762,  
13'd144,  -13'd374,  13'd182,  13'd294,  -13'd322,  -13'd744,  -13'd456,  13'd225,  -13'd674,  13'd257,  -13'd57,  -13'd198,  -13'd445,  13'd440,  13'd468,  -13'd571,  
-13'd384,  -13'd93,  -13'd329,  -13'd557,  13'd27,  -13'd413,  -13'd478,  13'd56,  -13'd596,  -13'd128,  13'd694,  -13'd295,  13'd281,  13'd903,  13'd197,  13'd404,  
13'd80,  -13'd823,  -13'd63,  13'd887,  13'd480,  13'd656,  -13'd376,  13'd448,  -13'd967,  -13'd156,  13'd246,  13'd140,  13'd621,  -13'd309,  13'd405,  13'd410,  
-13'd523,  13'd12,  -13'd76,  13'd257,  13'd754,  -13'd74,  13'd280,  13'd331,  13'd377,  13'd716,  13'd6,  13'd649,  13'd302,  -13'd180,  -13'd225,  -13'd78,  
13'd163,  13'd1168,  -13'd608,  13'd750,  13'd668,  13'd698,  13'd108,  -13'd25,  13'd789,  13'd901,  13'd276,  13'd126,  13'd98,  -13'd326,  13'd282,  13'd765,  

13'd136,  13'd291,  -13'd742,  -13'd152,  13'd112,  -13'd697,  -13'd514,  -13'd427,  13'd91,  -13'd34,  13'd129,  13'd445,  -13'd1083,  -13'd907,  -13'd563,  13'd2,  
13'd611,  -13'd488,  -13'd462,  13'd926,  -13'd151,  13'd95,  -13'd912,  13'd104,  -13'd217,  13'd229,  13'd487,  -13'd438,  13'd837,  -13'd343,  13'd8,  13'd664,  
-13'd315,  13'd257,  -13'd240,  13'd263,  -13'd12,  13'd737,  -13'd571,  13'd227,  13'd764,  13'd505,  -13'd681,  13'd397,  13'd558,  -13'd1697,  -13'd631,  13'd279,  
-13'd115,  -13'd58,  13'd73,  13'd117,  13'd507,  13'd102,  -13'd810,  13'd51,  -13'd548,  13'd633,  -13'd49,  13'd578,  13'd429,  -13'd729,  -13'd34,  -13'd629,  
-13'd1033,  -13'd471,  13'd839,  13'd211,  13'd558,  13'd30,  -13'd62,  13'd252,  -13'd412,  13'd438,  -13'd175,  -13'd140,  -13'd556,  -13'd38,  -13'd623,  -13'd739,  
13'd29,  -13'd467,  13'd319,  13'd679,  -13'd349,  13'd877,  13'd503,  13'd17,  13'd1155,  13'd439,  13'd175,  13'd312,  13'd380,  13'd12,  -13'd462,  -13'd341,  
-13'd305,  13'd1319,  -13'd337,  13'd26,  -13'd102,  -13'd524,  -13'd62,  13'd482,  13'd341,  -13'd22,  -13'd277,  13'd322,  13'd363,  -13'd149,  -13'd431,  13'd614,  
-13'd839,  13'd318,  13'd94,  -13'd502,  -13'd142,  13'd515,  -13'd138,  -13'd441,  -13'd423,  -13'd362,  13'd368,  13'd541,  13'd378,  -13'd224,  -13'd584,  13'd1250,  
13'd244,  13'd520,  13'd104,  -13'd466,  13'd241,  -13'd87,  13'd113,  -13'd245,  13'd668,  -13'd411,  13'd492,  13'd695,  -13'd277,  13'd639,  13'd394,  -13'd77,  
-13'd639,  -13'd344,  -13'd161,  13'd410,  -13'd80,  -13'd305,  13'd233,  -13'd315,  -13'd355,  -13'd632,  13'd30,  -13'd422,  -13'd371,  13'd19,  -13'd236,  13'd268,  
13'd676,  -13'd109,  13'd746,  13'd171,  13'd1253,  -13'd10,  13'd72,  13'd298,  13'd530,  13'd188,  -13'd105,  13'd208,  -13'd158,  -13'd243,  13'd293,  13'd418,  
-13'd80,  13'd444,  -13'd296,  -13'd231,  13'd378,  -13'd48,  13'd289,  13'd375,  -13'd1028,  -13'd291,  13'd688,  13'd234,  13'd41,  -13'd642,  13'd340,  -13'd633,  
13'd972,  -13'd207,  13'd900,  13'd280,  -13'd379,  -13'd201,  13'd248,  13'd132,  -13'd308,  13'd18,  13'd188,  -13'd348,  -13'd601,  13'd4,  13'd211,  -13'd695,  
13'd744,  13'd306,  13'd355,  -13'd660,  -13'd238,  -13'd193,  13'd763,  -13'd869,  13'd340,  -13'd707,  -13'd82,  13'd12,  -13'd62,  -13'd23,  -13'd519,  -13'd402,  
13'd1232,  13'd491,  13'd70,  -13'd305,  -13'd82,  13'd916,  13'd447,  -13'd115,  13'd290,  -13'd361,  13'd74,  13'd269,  -13'd272,  13'd898,  -13'd362,  13'd392,  
13'd93,  13'd394,  -13'd27,  13'd362,  13'd364,  -13'd624,  -13'd351,  13'd186,  -13'd427,  -13'd162,  13'd347,  13'd743,  13'd292,  13'd304,  13'd509,  -13'd610,  
-13'd90,  13'd904,  -13'd418,  -13'd454,  13'd453,  -13'd69,  -13'd313,  13'd465,  -13'd196,  -13'd1,  -13'd201,  13'd100,  -13'd563,  -13'd859,  13'd126,  13'd634,  
-13'd7,  13'd143,  -13'd620,  -13'd27,  13'd119,  -13'd419,  -13'd337,  13'd110,  13'd818,  13'd590,  -13'd619,  13'd478,  13'd143,  13'd425,  -13'd281,  13'd222,  
13'd682,  13'd254,  13'd6,  -13'd281,  -13'd157,  -13'd753,  13'd60,  -13'd332,  13'd677,  13'd430,  13'd324,  -13'd458,  -13'd408,  13'd2,  13'd112,  -13'd199,  
-13'd542,  -13'd719,  -13'd374,  -13'd117,  -13'd28,  -13'd1152,  13'd494,  -13'd225,  13'd645,  13'd198,  13'd502,  -13'd520,  13'd477,  13'd332,  -13'd509,  13'd332,  
13'd79,  -13'd74,  -13'd260,  -13'd229,  -13'd678,  -13'd88,  -13'd802,  -13'd675,  -13'd400,  13'd323,  13'd644,  -13'd194,  13'd168,  13'd692,  -13'd18,  -13'd52,  
13'd79,  -13'd40,  13'd345,  13'd103,  13'd652,  13'd94,  13'd189,  13'd26,  13'd267,  13'd264,  -13'd151,  13'd521,  -13'd206,  -13'd365,  13'd290,  13'd330,  
13'd307,  13'd92,  13'd542,  -13'd123,  -13'd28,  -13'd19,  13'd240,  13'd561,  13'd28,  -13'd575,  -13'd772,  -13'd623,  -13'd661,  -13'd34,  13'd45,  -13'd489,  
-13'd347,  -13'd244,  -13'd590,  -13'd390,  -13'd214,  13'd428,  -13'd46,  -13'd472,  13'd411,  -13'd335,  -13'd381,  13'd617,  13'd189,  13'd514,  13'd579,  -13'd414,  
-13'd214,  -13'd543,  13'd254,  13'd291,  -13'd240,  13'd126,  13'd68,  -13'd130,  -13'd759,  13'd902,  13'd193,  -13'd554,  13'd285,  13'd163,  13'd341,  -13'd73,  

-13'd122,  13'd442,  -13'd65,  13'd116,  -13'd643,  -13'd8,  13'd320,  -13'd49,  -13'd702,  -13'd109,  13'd1092,  13'd745,  13'd153,  13'd100,  13'd42,  13'd401,  
-13'd770,  13'd635,  -13'd336,  13'd40,  -13'd354,  -13'd3,  13'd240,  13'd29,  -13'd54,  13'd443,  13'd461,  13'd123,  -13'd191,  -13'd981,  13'd435,  -13'd10,  
-13'd21,  13'd464,  -13'd438,  -13'd617,  13'd980,  -13'd199,  13'd166,  13'd417,  13'd279,  13'd338,  13'd448,  -13'd149,  13'd135,  -13'd1444,  -13'd278,  -13'd158,  
-13'd484,  -13'd883,  13'd150,  13'd491,  -13'd58,  -13'd441,  -13'd332,  13'd587,  13'd53,  -13'd128,  -13'd83,  13'd508,  -13'd642,  13'd156,  -13'd257,  -13'd136,  
-13'd234,  -13'd640,  13'd502,  -13'd151,  -13'd630,  -13'd523,  -13'd96,  -13'd60,  -13'd39,  13'd134,  -13'd248,  13'd51,  -13'd22,  -13'd267,  -13'd175,  13'd585,  
13'd215,  13'd796,  -13'd380,  13'd75,  -13'd188,  13'd200,  -13'd705,  -13'd196,  -13'd62,  -13'd758,  13'd377,  -13'd7,  13'd676,  13'd535,  13'd427,  13'd848,  
13'd625,  13'd92,  -13'd383,  -13'd579,  13'd266,  -13'd68,  13'd364,  -13'd289,  13'd594,  -13'd745,  13'd274,  13'd428,  13'd55,  -13'd101,  13'd646,  13'd198,  
13'd561,  13'd424,  -13'd649,  13'd73,  13'd574,  -13'd229,  13'd197,  13'd555,  13'd499,  13'd224,  -13'd356,  13'd1157,  -13'd607,  -13'd171,  -13'd253,  13'd570,  
13'd224,  13'd238,  -13'd793,  -13'd135,  13'd286,  13'd106,  13'd860,  -13'd235,  -13'd75,  -13'd19,  -13'd514,  -13'd27,  13'd72,  -13'd193,  13'd116,  13'd177,  
-13'd769,  -13'd773,  -13'd419,  13'd226,  13'd179,  -13'd204,  13'd644,  -13'd19,  13'd228,  -13'd126,  -13'd41,  -13'd153,  13'd74,  13'd435,  -13'd656,  13'd94,  
-13'd336,  -13'd320,  13'd608,  13'd279,  -13'd201,  -13'd60,  13'd607,  -13'd408,  -13'd415,  -13'd176,  -13'd259,  -13'd500,  -13'd57,  -13'd48,  -13'd332,  -13'd583,  
13'd540,  -13'd139,  -13'd507,  13'd116,  -13'd110,  -13'd603,  -13'd591,  -13'd402,  -13'd582,  -13'd560,  -13'd26,  -13'd290,  13'd76,  13'd509,  13'd719,  13'd49,  
13'd361,  13'd2,  13'd352,  13'd94,  13'd246,  -13'd500,  -13'd116,  -13'd593,  -13'd208,  13'd34,  13'd493,  13'd165,  -13'd158,  13'd41,  -13'd283,  -13'd46,  
13'd520,  -13'd813,  -13'd221,  -13'd627,  13'd315,  13'd353,  -13'd608,  -13'd47,  13'd61,  -13'd21,  13'd293,  -13'd9,  -13'd126,  -13'd82,  13'd221,  13'd142,  
-13'd779,  -13'd67,  13'd366,  13'd218,  13'd462,  13'd482,  13'd6,  -13'd429,  -13'd5,  13'd685,  -13'd173,  13'd451,  -13'd346,  13'd15,  -13'd538,  -13'd23,  
13'd410,  13'd621,  13'd490,  13'd272,  13'd42,  -13'd23,  -13'd218,  -13'd297,  13'd649,  13'd436,  -13'd266,  -13'd1171,  13'd177,  -13'd236,  -13'd545,  -13'd216,  
-13'd506,  13'd73,  -13'd692,  -13'd257,  13'd615,  -13'd307,  13'd261,  13'd43,  -13'd141,  -13'd19,  13'd128,  -13'd188,  13'd210,  -13'd225,  -13'd778,  -13'd634,  
13'd95,  -13'd105,  13'd191,  -13'd299,  -13'd551,  -13'd525,  13'd96,  13'd750,  13'd112,  13'd40,  -13'd39,  -13'd517,  13'd413,  13'd549,  -13'd271,  13'd499,  
13'd679,  -13'd178,  13'd416,  13'd478,  13'd64,  13'd81,  -13'd676,  -13'd488,  -13'd328,  13'd195,  13'd432,  13'd600,  -13'd488,  13'd696,  13'd557,  13'd289,  
13'd504,  13'd713,  -13'd857,  13'd412,  -13'd203,  13'd241,  13'd326,  13'd663,  -13'd148,  13'd637,  -13'd97,  -13'd491,  13'd375,  13'd46,  13'd254,  -13'd318,  
13'd371,  13'd171,  -13'd446,  13'd56,  -13'd218,  -13'd491,  13'd248,  -13'd671,  13'd487,  -13'd156,  13'd420,  13'd1,  13'd41,  -13'd993,  13'd360,  13'd384,  
13'd561,  13'd654,  13'd133,  -13'd544,  -13'd885,  -13'd393,  13'd393,  -13'd921,  13'd1136,  -13'd463,  -13'd714,  -13'd172,  -13'd331,  -13'd584,  -13'd676,  13'd347,  
-13'd574,  13'd229,  13'd520,  -13'd421,  -13'd259,  13'd238,  13'd14,  -13'd152,  13'd1044,  13'd1405,  -13'd741,  13'd299,  13'd15,  13'd1303,  13'd438,  -13'd81,  
13'd513,  -13'd503,  13'd187,  -13'd53,  -13'd170,  13'd20,  13'd392,  13'd560,  13'd709,  -13'd400,  -13'd485,  13'd699,  -13'd24,  13'd792,  -13'd583,  -13'd329,  
-13'd392,  13'd660,  13'd899,  13'd709,  13'd191,  -13'd203,  13'd828,  13'd703,  13'd699,  -13'd180,  -13'd679,  -13'd55,  13'd413,  13'd170,  13'd187,  13'd66,  

-13'd412,  -13'd289,  -13'd419,  13'd325,  13'd486,  -13'd309,  -13'd1446,  13'd223,  -13'd381,  -13'd131,  -13'd539,  -13'd62,  13'd331,  -13'd194,  13'd720,  13'd543,  
-13'd359,  -13'd181,  -13'd165,  13'd170,  -13'd293,  -13'd475,  -13'd45,  13'd797,  -13'd166,  13'd739,  -13'd229,  -13'd156,  13'd155,  -13'd849,  -13'd256,  -13'd46,  
-13'd424,  13'd484,  13'd277,  13'd969,  13'd55,  -13'd470,  -13'd634,  13'd763,  -13'd503,  -13'd331,  -13'd721,  13'd210,  13'd199,  -13'd1233,  -13'd83,  13'd726,  
13'd250,  -13'd304,  -13'd319,  13'd473,  -13'd232,  13'd496,  -13'd275,  13'd269,  -13'd30,  13'd420,  13'd500,  13'd166,  13'd580,  -13'd600,  -13'd88,  13'd1142,  
-13'd168,  -13'd870,  13'd166,  13'd48,  13'd24,  13'd84,  13'd601,  -13'd436,  13'd418,  13'd1070,  13'd167,  13'd341,  13'd349,  -13'd244,  -13'd198,  13'd99,  
-13'd521,  13'd303,  13'd48,  13'd502,  13'd558,  13'd58,  -13'd699,  -13'd500,  13'd325,  13'd233,  -13'd409,  13'd768,  13'd673,  -13'd748,  -13'd920,  13'd482,  
-13'd294,  -13'd68,  -13'd248,  -13'd177,  13'd263,  13'd42,  13'd315,  -13'd41,  -13'd26,  -13'd470,  13'd193,  -13'd398,  13'd435,  -13'd726,  -13'd676,  13'd206,  
-13'd12,  13'd126,  -13'd398,  13'd340,  13'd142,  -13'd74,  13'd281,  -13'd180,  -13'd826,  13'd729,  13'd354,  -13'd379,  13'd355,  13'd1043,  13'd50,  13'd411,  
13'd103,  13'd168,  13'd1054,  -13'd425,  -13'd60,  13'd523,  13'd207,  -13'd180,  -13'd372,  13'd142,  13'd144,  13'd541,  13'd58,  13'd348,  13'd481,  13'd1155,  
13'd2,  -13'd78,  -13'd511,  13'd385,  13'd12,  13'd338,  13'd686,  13'd390,  13'd54,  -13'd203,  -13'd207,  13'd23,  -13'd28,  13'd416,  13'd132,  -13'd232,  
-13'd545,  13'd543,  -13'd655,  13'd215,  -13'd148,  -13'd110,  13'd62,  13'd421,  13'd856,  -13'd784,  13'd140,  13'd65,  -13'd301,  -13'd724,  -13'd493,  13'd277,  
13'd156,  -13'd730,  -13'd334,  -13'd1032,  13'd768,  13'd0,  13'd131,  -13'd141,  13'd95,  -13'd228,  -13'd13,  -13'd315,  13'd604,  -13'd130,  13'd261,  13'd138,  
-13'd276,  -13'd365,  13'd690,  13'd324,  13'd386,  13'd19,  -13'd318,  -13'd767,  -13'd364,  -13'd128,  -13'd603,  13'd22,  -13'd419,  13'd392,  13'd393,  -13'd309,  
13'd406,  13'd636,  13'd244,  -13'd315,  13'd814,  13'd687,  13'd367,  13'd728,  13'd466,  13'd583,  13'd111,  13'd358,  13'd647,  13'd210,  -13'd138,  13'd10,  
13'd846,  -13'd204,  13'd748,  -13'd2,  13'd411,  13'd553,  13'd521,  13'd153,  -13'd626,  -13'd591,  -13'd126,  13'd542,  13'd469,  13'd30,  13'd448,  13'd277,  
13'd179,  13'd74,  -13'd80,  13'd431,  -13'd449,  -13'd239,  13'd214,  13'd359,  13'd293,  13'd176,  -13'd392,  13'd277,  -13'd603,  -13'd241,  13'd229,  13'd109,  
13'd715,  13'd20,  -13'd19,  -13'd296,  -13'd185,  13'd319,  -13'd489,  13'd7,  13'd392,  13'd206,  13'd137,  -13'd200,  13'd9,  13'd306,  -13'd2,  -13'd371,  
-13'd346,  13'd123,  13'd303,  13'd557,  13'd39,  -13'd542,  13'd73,  13'd579,  13'd71,  -13'd696,  13'd574,  -13'd193,  -13'd113,  -13'd169,  -13'd16,  -13'd218,  
-13'd737,  -13'd628,  13'd62,  13'd49,  -13'd288,  -13'd339,  13'd522,  -13'd258,  -13'd504,  -13'd555,  13'd789,  13'd483,  13'd417,  13'd21,  13'd634,  -13'd137,  
13'd318,  -13'd81,  -13'd140,  -13'd787,  13'd265,  13'd126,  13'd403,  -13'd324,  -13'd679,  -13'd195,  13'd580,  -13'd49,  -13'd70,  -13'd533,  -13'd239,  13'd325,  
-13'd172,  13'd77,  -13'd16,  -13'd179,  13'd7,  -13'd370,  -13'd237,  -13'd35,  -13'd628,  13'd14,  -13'd63,  -13'd74,  -13'd447,  -13'd468,  13'd670,  13'd215,  
-13'd175,  13'd246,  -13'd263,  -13'd122,  -13'd136,  -13'd720,  -13'd18,  -13'd786,  13'd300,  -13'd684,  -13'd109,  13'd195,  13'd385,  13'd191,  -13'd562,  13'd486,  
13'd63,  13'd248,  13'd237,  -13'd757,  -13'd679,  -13'd789,  -13'd92,  13'd401,  -13'd42,  13'd839,  -13'd815,  13'd373,  -13'd540,  13'd211,  -13'd662,  -13'd26,  
-13'd331,  13'd310,  13'd404,  -13'd329,  13'd323,  -13'd101,  13'd430,  -13'd254,  -13'd625,  -13'd114,  13'd35,  13'd200,  -13'd582,  -13'd605,  13'd242,  -13'd514,  
13'd206,  13'd412,  13'd6,  -13'd796,  13'd15,  -13'd886,  -13'd283,  -13'd112,  -13'd600,  -13'd342,  13'd273,  -13'd1134,  -13'd457,  -13'd312,  -13'd877,  -13'd179,  

-13'd414,  13'd582,  -13'd109,  13'd154,  13'd413,  13'd427,  -13'd394,  -13'd45,  13'd754,  13'd165,  13'd130,  -13'd577,  -13'd144,  13'd312,  -13'd249,  -13'd383,  
-13'd529,  -13'd211,  13'd893,  13'd663,  13'd288,  13'd235,  13'd293,  13'd43,  -13'd196,  -13'd201,  -13'd333,  13'd8,  13'd788,  13'd197,  13'd759,  13'd758,  
13'd379,  -13'd635,  13'd459,  -13'd410,  -13'd56,  13'd241,  13'd757,  13'd215,  13'd247,  13'd642,  13'd474,  13'd449,  -13'd183,  13'd706,  13'd549,  -13'd390,  
13'd398,  -13'd226,  -13'd151,  13'd617,  -13'd362,  -13'd103,  13'd271,  -13'd560,  13'd888,  13'd90,  13'd257,  -13'd453,  -13'd167,  13'd789,  -13'd1040,  -13'd279,  
13'd215,  -13'd165,  -13'd573,  -13'd768,  13'd529,  -13'd574,  13'd746,  13'd134,  13'd30,  -13'd334,  13'd496,  -13'd204,  13'd289,  -13'd354,  -13'd500,  -13'd284,  
-13'd728,  -13'd395,  -13'd234,  -13'd854,  13'd683,  -13'd538,  13'd203,  13'd416,  -13'd428,  13'd180,  13'd150,  -13'd853,  -13'd467,  -13'd608,  13'd75,  13'd58,  
-13'd376,  -13'd359,  13'd79,  13'd254,  -13'd152,  -13'd440,  -13'd1365,  -13'd256,  -13'd635,  13'd604,  -13'd306,  -13'd651,  -13'd347,  -13'd1095,  13'd23,  13'd16,  
13'd454,  -13'd1295,  13'd796,  13'd249,  -13'd43,  13'd711,  13'd65,  13'd16,  -13'd1555,  13'd43,  13'd90,  -13'd183,  -13'd314,  13'd182,  13'd393,  13'd177,  
13'd864,  -13'd401,  13'd698,  13'd407,  13'd85,  -13'd333,  13'd546,  13'd1068,  -13'd872,  -13'd145,  13'd478,  -13'd579,  -13'd303,  13'd577,  13'd69,  -13'd59,  
13'd1220,  -13'd524,  13'd433,  13'd538,  -13'd303,  -13'd62,  -13'd342,  -13'd160,  13'd406,  13'd458,  13'd290,  -13'd632,  -13'd135,  13'd201,  -13'd678,  -13'd14,  
-13'd727,  -13'd259,  -13'd1013,  -13'd4,  13'd402,  -13'd587,  -13'd240,  13'd242,  13'd500,  13'd80,  -13'd149,  -13'd1234,  13'd146,  -13'd1298,  -13'd331,  -13'd590,  
-13'd47,  -13'd352,  -13'd278,  13'd244,  -13'd810,  13'd69,  -13'd810,  -13'd255,  13'd149,  13'd171,  13'd102,  13'd151,  -13'd809,  -13'd72,  13'd381,  13'd331,  
13'd917,  13'd391,  13'd635,  13'd112,  -13'd869,  13'd17,  -13'd784,  13'd256,  -13'd257,  13'd833,  13'd501,  -13'd230,  13'd261,  -13'd106,  13'd1017,  13'd381,  
13'd349,  -13'd444,  13'd156,  13'd133,  -13'd114,  13'd87,  -13'd340,  13'd445,  -13'd542,  13'd545,  -13'd282,  -13'd648,  13'd998,  -13'd517,  -13'd418,  13'd244,  
-13'd513,  -13'd380,  -13'd49,  13'd385,  -13'd591,  -13'd563,  13'd323,  13'd258,  13'd543,  -13'd130,  13'd436,  -13'd98,  -13'd124,  13'd81,  -13'd315,  -13'd17,  
-13'd1019,  -13'd45,  -13'd507,  13'd179,  13'd99,  13'd205,  13'd54,  13'd287,  13'd266,  13'd461,  13'd313,  -13'd892,  -13'd662,  13'd389,  13'd133,  -13'd327,  
13'd371,  13'd499,  -13'd253,  -13'd108,  -13'd468,  13'd613,  13'd197,  -13'd49,  -13'd528,  13'd230,  13'd145,  -13'd88,  13'd226,  -13'd111,  13'd217,  -13'd296,  
13'd306,  -13'd14,  -13'd594,  13'd355,  -13'd278,  -13'd35,  13'd249,  13'd366,  -13'd84,  13'd175,  13'd322,  13'd112,  13'd612,  -13'd752,  13'd216,  13'd338,  
-13'd7,  -13'd298,  13'd759,  13'd203,  -13'd491,  -13'd308,  -13'd458,  -13'd186,  -13'd366,  13'd115,  13'd462,  13'd64,  -13'd377,  -13'd106,  13'd14,  13'd20,  
-13'd408,  -13'd135,  13'd5,  -13'd118,  13'd150,  -13'd208,  13'd120,  13'd544,  -13'd372,  13'd637,  -13'd63,  -13'd200,  -13'd48,  13'd341,  -13'd383,  -13'd125,  
13'd212,  13'd738,  -13'd222,  13'd440,  -13'd102,  13'd383,  13'd519,  -13'd225,  13'd467,  -13'd129,  -13'd351,  13'd632,  13'd166,  -13'd274,  13'd218,  -13'd85,  
13'd28,  13'd530,  13'd170,  -13'd63,  13'd170,  -13'd42,  13'd253,  13'd205,  -13'd297,  -13'd137,  -13'd547,  13'd54,  13'd173,  13'd474,  13'd502,  -13'd326,  
13'd357,  -13'd208,  13'd244,  -13'd338,  13'd357,  13'd295,  13'd263,  -13'd277,  13'd351,  13'd550,  13'd381,  -13'd81,  -13'd324,  -13'd445,  13'd417,  13'd360,  
-13'd234,  13'd270,  -13'd41,  -13'd376,  -13'd476,  -13'd807,  13'd526,  -13'd511,  -13'd475,  -13'd337,  13'd142,  13'd120,  -13'd451,  13'd881,  13'd264,  13'd276,  
13'd319,  13'd706,  -13'd40,  13'd354,  13'd257,  -13'd669,  -13'd438,  -13'd294,  13'd738,  -13'd416,  13'd264,  -13'd127,  -13'd913,  13'd641,  -13'd452,  -13'd46,  

-13'd669,  13'd415,  -13'd285,  -13'd406,  -13'd196,  13'd1,  -13'd173,  -13'd659,  -13'd463,  -13'd702,  -13'd1065,  -13'd499,  -13'd340,  -13'd648,  -13'd435,  -13'd439,  
-13'd561,  13'd466,  -13'd126,  13'd548,  -13'd134,  13'd820,  13'd190,  13'd172,  13'd357,  -13'd130,  -13'd1183,  13'd137,  -13'd526,  13'd252,  13'd58,  13'd202,  
13'd467,  -13'd66,  -13'd254,  13'd87,  13'd912,  13'd645,  13'd497,  -13'd576,  -13'd779,  -13'd478,  13'd465,  13'd346,  -13'd559,  -13'd365,  13'd374,  -13'd740,  
-13'd455,  -13'd195,  -13'd38,  13'd603,  -13'd48,  13'd618,  -13'd383,  -13'd115,  -13'd171,  -13'd228,  13'd342,  -13'd314,  13'd769,  13'd1263,  -13'd328,  -13'd668,  
-13'd458,  -13'd735,  -13'd218,  13'd578,  13'd722,  -13'd158,  13'd225,  13'd41,  -13'd702,  13'd363,  -13'd305,  -13'd686,  -13'd389,  -13'd198,  13'd303,  -13'd787,  
-13'd462,  -13'd276,  -13'd831,  13'd151,  13'd862,  -13'd854,  -13'd177,  -13'd809,  13'd161,  -13'd244,  -13'd66,  13'd343,  -13'd188,  -13'd60,  -13'd746,  -13'd877,  
13'd407,  -13'd108,  13'd351,  -13'd809,  13'd550,  -13'd305,  -13'd208,  -13'd356,  -13'd482,  13'd221,  -13'd572,  -13'd894,  -13'd963,  -13'd505,  -13'd207,  -13'd795,  
13'd346,  13'd628,  13'd424,  13'd20,  -13'd937,  13'd72,  -13'd89,  13'd247,  13'd462,  13'd337,  -13'd188,  -13'd387,  -13'd294,  13'd315,  13'd465,  -13'd620,  
13'd27,  13'd13,  13'd558,  13'd147,  -13'd102,  -13'd358,  13'd637,  -13'd288,  -13'd315,  -13'd294,  13'd446,  13'd605,  13'd197,  13'd1234,  13'd376,  13'd369,  
-13'd349,  13'd254,  13'd301,  -13'd276,  -13'd17,  -13'd186,  13'd311,  -13'd579,  13'd184,  -13'd170,  -13'd44,  13'd120,  -13'd286,  -13'd123,  -13'd652,  -13'd514,  
-13'd687,  -13'd593,  -13'd17,  13'd321,  13'd76,  -13'd321,  -13'd69,  13'd115,  13'd702,  -13'd294,  13'd249,  -13'd220,  -13'd143,  13'd312,  -13'd71,  -13'd662,  
-13'd169,  -13'd554,  13'd49,  13'd451,  13'd344,  13'd762,  13'd161,  -13'd133,  13'd447,  -13'd133,  -13'd148,  -13'd404,  13'd118,  -13'd315,  13'd182,  13'd230,  
13'd458,  13'd55,  13'd402,  -13'd394,  13'd327,  13'd808,  -13'd40,  13'd562,  13'd594,  -13'd117,  -13'd586,  13'd448,  -13'd0,  13'd125,  13'd415,  -13'd641,  
13'd288,  -13'd250,  13'd242,  -13'd88,  -13'd12,  13'd264,  13'd327,  13'd281,  13'd579,  13'd105,  -13'd365,  -13'd47,  13'd481,  13'd520,  13'd289,  -13'd391,  
13'd419,  13'd637,  -13'd67,  13'd238,  13'd111,  -13'd953,  -13'd388,  -13'd16,  -13'd713,  -13'd995,  13'd134,  -13'd457,  -13'd265,  -13'd404,  -13'd17,  13'd62,  
13'd397,  -13'd190,  13'd416,  13'd129,  -13'd296,  -13'd491,  13'd570,  -13'd561,  13'd157,  -13'd984,  13'd1134,  13'd628,  13'd237,  -13'd253,  -13'd168,  13'd324,  
13'd224,  -13'd192,  -13'd7,  -13'd473,  -13'd1217,  13'd113,  13'd556,  -13'd52,  13'd204,  13'd177,  13'd535,  -13'd595,  13'd419,  13'd619,  13'd197,  13'd796,  
13'd393,  -13'd405,  -13'd431,  13'd479,  -13'd423,  13'd584,  13'd138,  13'd908,  13'd554,  -13'd391,  13'd569,  -13'd455,  13'd242,  13'd600,  13'd648,  13'd193,  
-13'd171,  -13'd376,  -13'd468,  -13'd25,  -13'd182,  13'd116,  13'd354,  13'd695,  -13'd371,  13'd473,  -13'd37,  13'd68,  -13'd156,  13'd688,  -13'd168,  -13'd127,  
13'd556,  13'd319,  -13'd192,  13'd162,  -13'd1230,  -13'd364,  -13'd1039,  -13'd630,  -13'd1063,  -13'd1156,  13'd216,  13'd327,  -13'd828,  13'd859,  -13'd207,  -13'd387,  
13'd134,  -13'd934,  13'd86,  -13'd546,  -13'd606,  13'd134,  13'd779,  -13'd276,  13'd138,  13'd194,  13'd254,  -13'd3,  -13'd445,  13'd473,  13'd10,  -13'd379,  
13'd450,  13'd195,  -13'd44,  -13'd674,  13'd171,  13'd235,  13'd861,  -13'd712,  13'd989,  13'd750,  13'd23,  -13'd79,  -13'd657,  13'd8,  -13'd255,  13'd173,  
13'd62,  -13'd264,  13'd1079,  -13'd641,  13'd437,  -13'd304,  -13'd130,  13'd325,  13'd509,  13'd498,  -13'd610,  13'd102,  -13'd509,  13'd552,  13'd430,  -13'd501,  
-13'd1152,  -13'd591,  -13'd210,  13'd393,  13'd723,  -13'd190,  13'd612,  -13'd76,  13'd44,  13'd212,  -13'd340,  -13'd615,  13'd49,  -13'd165,  13'd74,  -13'd515,  
13'd5,  13'd258,  13'd831,  13'd213,  -13'd12,  13'd184,  -13'd412,  13'd124,  13'd37,  13'd354,  -13'd626,  13'd271,  13'd787,  13'd82,  -13'd398,  13'd111,  

-13'd458,  -13'd213,  -13'd593,  13'd630,  13'd539,  -13'd364,  13'd176,  13'd407,  -13'd666,  -13'd489,  13'd740,  -13'd973,  13'd265,  -13'd619,  -13'd426,  13'd20,  
13'd112,  -13'd269,  -13'd417,  13'd600,  13'd165,  13'd417,  -13'd189,  13'd276,  13'd92,  -13'd274,  -13'd643,  -13'd34,  13'd672,  -13'd1051,  -13'd278,  -13'd437,  
-13'd391,  -13'd532,  -13'd629,  13'd279,  -13'd7,  -13'd244,  -13'd791,  -13'd49,  -13'd471,  -13'd299,  13'd341,  -13'd802,  -13'd253,  -13'd649,  -13'd435,  13'd232,  
-13'd431,  -13'd1065,  13'd502,  13'd516,  13'd392,  -13'd11,  13'd129,  -13'd297,  -13'd287,  13'd643,  13'd201,  -13'd95,  -13'd240,  -13'd401,  13'd664,  13'd482,  
-13'd452,  -13'd875,  13'd310,  -13'd112,  -13'd123,  -13'd90,  -13'd57,  -13'd510,  13'd554,  -13'd489,  -13'd106,  -13'd10,  -13'd771,  13'd28,  -13'd18,  -13'd118,  
-13'd431,  13'd96,  -13'd908,  13'd15,  -13'd625,  -13'd808,  13'd21,  -13'd329,  -13'd103,  -13'd235,  13'd974,  -13'd323,  13'd217,  13'd63,  -13'd413,  -13'd725,  
-13'd197,  -13'd621,  -13'd284,  13'd192,  13'd387,  -13'd768,  13'd322,  -13'd624,  -13'd176,  13'd287,  -13'd189,  13'd872,  -13'd406,  -13'd855,  13'd452,  13'd181,  
-13'd87,  13'd275,  -13'd195,  13'd82,  13'd722,  13'd299,  13'd238,  -13'd104,  13'd173,  13'd438,  13'd216,  13'd699,  13'd434,  13'd22,  13'd194,  13'd468,  
13'd509,  -13'd439,  -13'd689,  -13'd171,  13'd862,  13'd138,  -13'd26,  13'd462,  -13'd126,  13'd479,  13'd3,  13'd905,  13'd56,  13'd92,  -13'd58,  13'd99,  
-13'd572,  13'd535,  13'd583,  13'd811,  -13'd39,  13'd83,  13'd843,  13'd151,  13'd260,  13'd769,  13'd149,  13'd604,  -13'd146,  -13'd226,  13'd627,  13'd101,  
-13'd430,  13'd460,  13'd585,  13'd402,  -13'd415,  13'd83,  -13'd414,  -13'd329,  13'd124,  -13'd337,  13'd109,  -13'd242,  -13'd474,  -13'd741,  -13'd644,  -13'd497,  
13'd13,  -13'd62,  -13'd88,  -13'd301,  -13'd338,  -13'd92,  -13'd713,  13'd123,  -13'd57,  13'd206,  -13'd678,  13'd191,  -13'd508,  -13'd1113,  -13'd243,  -13'd89,  
13'd799,  -13'd774,  -13'd262,  -13'd422,  -13'd247,  -13'd950,  -13'd393,  -13'd13,  13'd178,  13'd381,  13'd179,  -13'd128,  -13'd154,  -13'd421,  13'd628,  13'd477,  
-13'd312,  -13'd120,  13'd246,  -13'd441,  13'd443,  13'd250,  13'd91,  13'd518,  -13'd477,  13'd89,  13'd497,  -13'd134,  13'd239,  -13'd442,  -13'd36,  13'd307,  
-13'd78,  -13'd361,  -13'd19,  13'd540,  13'd567,  13'd45,  -13'd218,  13'd584,  13'd47,  13'd15,  -13'd168,  13'd530,  -13'd447,  13'd81,  13'd0,  -13'd34,  
-13'd422,  -13'd318,  13'd95,  -13'd41,  -13'd522,  13'd520,  -13'd1022,  13'd380,  13'd589,  13'd26,  -13'd341,  -13'd548,  13'd696,  13'd518,  -13'd525,  13'd189,  
-13'd119,  -13'd956,  -13'd719,  13'd265,  -13'd23,  -13'd321,  -13'd545,  13'd667,  -13'd666,  13'd431,  13'd535,  13'd293,  13'd341,  -13'd113,  -13'd32,  13'd331,  
-13'd719,  13'd269,  -13'd276,  -13'd326,  13'd511,  -13'd649,  -13'd63,  13'd369,  -13'd374,  -13'd474,  13'd69,  -13'd380,  13'd387,  -13'd426,  13'd511,  -13'd450,  
13'd297,  13'd410,  13'd340,  13'd48,  13'd668,  13'd265,  -13'd248,  -13'd227,  -13'd210,  13'd426,  -13'd217,  13'd191,  -13'd296,  13'd102,  13'd269,  13'd305,  
13'd111,  -13'd135,  13'd477,  -13'd312,  -13'd47,  -13'd160,  13'd458,  13'd21,  -13'd354,  13'd577,  13'd475,  -13'd407,  13'd778,  -13'd215,  13'd282,  -13'd83,  
-13'd381,  -13'd35,  13'd229,  -13'd118,  13'd20,  13'd223,  -13'd569,  13'd153,  13'd142,  13'd224,  -13'd48,  -13'd203,  13'd288,  13'd112,  13'd583,  -13'd224,  
13'd5,  13'd59,  13'd55,  13'd397,  13'd453,  -13'd60,  13'd605,  -13'd522,  -13'd894,  -13'd537,  -13'd11,  13'd676,  13'd157,  -13'd578,  -13'd367,  13'd1,  
-13'd65,  13'd70,  13'd100,  13'd83,  13'd602,  13'd178,  -13'd36,  -13'd552,  -13'd91,  13'd327,  -13'd247,  13'd802,  13'd711,  -13'd446,  -13'd46,  13'd594,  
13'd479,  13'd770,  -13'd380,  -13'd347,  13'd286,  13'd198,  13'd126,  -13'd652,  13'd500,  -13'd23,  -13'd95,  -13'd394,  13'd394,  -13'd204,  -13'd362,  13'd637,  
13'd775,  13'd1183,  13'd421,  -13'd84,  13'd573,  13'd502,  -13'd130,  13'd657,  13'd1063,  13'd1502,  -13'd309,  13'd742,  -13'd662,  13'd794,  13'd215,  13'd403,  

13'd168,  13'd144,  13'd884,  13'd168,  -13'd127,  13'd150,  13'd412,  -13'd200,  13'd316,  13'd471,  -13'd194,  -13'd179,  13'd161,  13'd268,  -13'd622,  13'd355,  
-13'd61,  -13'd160,  13'd203,  -13'd308,  -13'd392,  13'd14,  13'd252,  -13'd243,  -13'd375,  -13'd104,  13'd722,  13'd17,  -13'd337,  13'd1247,  -13'd772,  13'd107,  
-13'd257,  -13'd934,  13'd562,  -13'd207,  -13'd871,  -13'd214,  13'd469,  13'd403,  -13'd188,  13'd449,  13'd612,  -13'd448,  13'd703,  13'd808,  -13'd433,  -13'd708,  
13'd687,  13'd844,  -13'd281,  13'd67,  13'd199,  -13'd272,  13'd366,  13'd358,  -13'd5,  -13'd136,  13'd558,  13'd739,  13'd45,  -13'd85,  -13'd378,  -13'd205,  
13'd1400,  13'd1028,  -13'd438,  13'd401,  -13'd256,  13'd785,  -13'd98,  13'd182,  -13'd534,  13'd133,  -13'd29,  13'd693,  13'd459,  13'd155,  13'd301,  13'd77,  
13'd103,  13'd42,  13'd63,  13'd294,  -13'd302,  13'd663,  13'd731,  13'd17,  13'd149,  -13'd144,  13'd65,  13'd11,  -13'd111,  13'd492,  13'd710,  -13'd211,  
13'd202,  -13'd762,  -13'd208,  13'd340,  -13'd2,  13'd331,  13'd383,  13'd274,  13'd149,  -13'd442,  13'd1061,  13'd33,  -13'd306,  13'd42,  13'd433,  -13'd694,  
-13'd584,  -13'd226,  -13'd230,  -13'd174,  -13'd1080,  -13'd17,  -13'd169,  -13'd680,  13'd252,  13'd36,  13'd374,  -13'd1023,  13'd439,  13'd251,  -13'd254,  -13'd534,  
-13'd111,  -13'd132,  -13'd883,  13'd406,  13'd309,  -13'd686,  -13'd359,  13'd231,  -13'd15,  13'd151,  13'd280,  13'd96,  13'd290,  -13'd13,  -13'd344,  -13'd327,  
13'd180,  -13'd948,  -13'd622,  13'd251,  13'd44,  13'd576,  -13'd807,  -13'd423,  13'd301,  13'd147,  -13'd185,  13'd402,  -13'd44,  -13'd119,  -13'd527,  13'd936,  
-13'd413,  13'd304,  13'd248,  13'd457,  -13'd5,  13'd345,  13'd237,  13'd296,  -13'd506,  -13'd471,  -13'd31,  13'd145,  13'd756,  13'd418,  13'd767,  13'd179,  
13'd280,  -13'd515,  13'd130,  13'd100,  13'd673,  13'd104,  -13'd62,  13'd594,  13'd166,  -13'd335,  13'd1038,  13'd246,  -13'd68,  -13'd604,  -13'd92,  13'd324,  
-13'd287,  -13'd240,  -13'd457,  13'd441,  -13'd256,  -13'd675,  13'd4,  -13'd207,  -13'd258,  13'd693,  13'd322,  -13'd153,  -13'd402,  13'd32,  -13'd943,  -13'd104,  
-13'd373,  13'd90,  -13'd454,  13'd546,  13'd866,  13'd142,  13'd140,  -13'd325,  13'd79,  13'd451,  13'd230,  13'd39,  -13'd284,  13'd407,  13'd410,  13'd7,  
-13'd745,  -13'd151,  13'd338,  13'd600,  -13'd70,  -13'd628,  -13'd676,  -13'd318,  13'd256,  13'd823,  13'd89,  -13'd516,  -13'd477,  -13'd158,  13'd221,  13'd161,  
-13'd209,  13'd383,  -13'd416,  13'd549,  13'd512,  -13'd300,  13'd145,  13'd644,  13'd53,  -13'd31,  -13'd7,  -13'd866,  13'd630,  -13'd106,  -13'd117,  13'd929,  
-13'd929,  13'd816,  -13'd161,  13'd354,  13'd319,  -13'd106,  13'd29,  -13'd3,  -13'd192,  -13'd561,  -13'd863,  13'd537,  13'd355,  -13'd747,  -13'd410,  13'd143,  
-13'd587,  -13'd290,  -13'd590,  -13'd366,  13'd507,  13'd381,  -13'd144,  -13'd148,  13'd115,  13'd401,  13'd220,  13'd722,  13'd389,  13'd810,  -13'd21,  13'd726,  
13'd91,  -13'd763,  13'd61,  -13'd275,  13'd582,  13'd2,  13'd175,  13'd91,  13'd322,  13'd87,  13'd450,  13'd725,  13'd153,  13'd62,  -13'd180,  13'd721,  
-13'd461,  13'd2,  13'd782,  -13'd276,  13'd568,  13'd45,  13'd722,  -13'd50,  13'd59,  13'd337,  13'd92,  -13'd296,  -13'd318,  13'd154,  -13'd391,  13'd128,  
13'd399,  -13'd211,  -13'd665,  -13'd721,  13'd303,  -13'd193,  13'd613,  -13'd349,  13'd363,  13'd155,  13'd153,  13'd488,  -13'd342,  -13'd966,  -13'd324,  13'd167,  
13'd224,  13'd621,  -13'd188,  -13'd619,  13'd783,  13'd231,  13'd792,  13'd318,  13'd165,  -13'd439,  -13'd456,  -13'd135,  13'd178,  -13'd276,  -13'd180,  13'd112,  
-13'd306,  13'd75,  13'd337,  -13'd172,  13'd555,  -13'd875,  13'd475,  -13'd233,  13'd410,  13'd414,  -13'd234,  13'd294,  13'd116,  13'd59,  13'd594,  13'd74,  
13'd566,  -13'd167,  13'd762,  -13'd49,  13'd37,  -13'd657,  -13'd308,  13'd92,  -13'd52,  13'd516,  13'd382,  -13'd371,  13'd380,  13'd939,  -13'd209,  -13'd95,  
13'd579,  -13'd89,  -13'd338,  -13'd161,  -13'd191,  13'd930,  13'd96,  13'd390,  -13'd99,  -13'd22,  -13'd340,  13'd253,  -13'd322,  13'd438,  13'd943,  -13'd261,  

-13'd827,  -13'd920,  -13'd324,  -13'd314,  13'd249,  -13'd226,  -13'd765,  -13'd189,  13'd157,  13'd188,  -13'd701,  -13'd401,  -13'd1021,  -13'd759,  13'd258,  -13'd113,  
13'd359,  -13'd176,  13'd325,  -13'd260,  -13'd122,  13'd577,  13'd60,  -13'd104,  -13'd410,  -13'd99,  -13'd656,  13'd742,  13'd412,  13'd540,  -13'd500,  -13'd38,  
13'd451,  -13'd332,  13'd308,  13'd334,  13'd236,  -13'd166,  -13'd146,  -13'd354,  13'd59,  -13'd687,  -13'd347,  13'd642,  -13'd8,  -13'd66,  -13'd51,  -13'd582,  
13'd690,  -13'd816,  -13'd418,  13'd56,  -13'd147,  13'd101,  13'd760,  -13'd170,  -13'd74,  13'd752,  13'd53,  13'd75,  13'd25,  13'd1442,  13'd116,  -13'd715,  
-13'd917,  13'd510,  13'd513,  -13'd76,  13'd175,  -13'd336,  -13'd461,  13'd17,  13'd46,  13'd517,  13'd134,  -13'd398,  -13'd788,  -13'd129,  13'd164,  -13'd614,  
13'd401,  13'd583,  -13'd149,  -13'd138,  13'd318,  13'd583,  13'd345,  -13'd896,  13'd706,  -13'd232,  13'd334,  13'd530,  -13'd891,  13'd315,  -13'd276,  13'd62,  
-13'd294,  13'd656,  13'd371,  -13'd277,  -13'd447,  13'd768,  -13'd542,  13'd431,  -13'd374,  13'd708,  -13'd610,  13'd133,  13'd484,  13'd322,  -13'd122,  -13'd374,  
13'd670,  -13'd687,  13'd350,  13'd19,  -13'd419,  13'd785,  13'd571,  13'd478,  -13'd888,  13'd55,  -13'd183,  13'd536,  -13'd488,  -13'd89,  -13'd27,  -13'd247,  
13'd527,  13'd402,  13'd986,  13'd267,  13'd649,  13'd18,  13'd573,  13'd62,  -13'd377,  -13'd518,  13'd22,  13'd173,  13'd136,  13'd521,  -13'd222,  -13'd263,  
13'd361,  13'd202,  13'd802,  13'd324,  -13'd192,  -13'd339,  13'd45,  13'd423,  -13'd385,  -13'd826,  13'd334,  13'd328,  13'd57,  13'd269,  13'd72,  -13'd841,  
13'd121,  -13'd150,  13'd69,  -13'd37,  13'd717,  -13'd808,  13'd371,  -13'd175,  -13'd211,  -13'd378,  -13'd396,  -13'd63,  -13'd296,  -13'd9,  13'd525,  13'd295,  
13'd880,  13'd171,  13'd857,  13'd132,  13'd276,  -13'd571,  13'd520,  -13'd149,  -13'd124,  -13'd118,  13'd73,  13'd108,  13'd141,  13'd700,  13'd813,  -13'd37,  
13'd610,  13'd371,  13'd462,  13'd4,  -13'd785,  13'd483,  -13'd119,  13'd238,  -13'd180,  13'd272,  -13'd241,  -13'd203,  -13'd189,  13'd258,  13'd298,  -13'd298,  
-13'd91,  -13'd386,  13'd1018,  13'd559,  -13'd185,  -13'd335,  13'd206,  13'd376,  -13'd336,  13'd569,  13'd313,  -13'd782,  -13'd108,  13'd454,  13'd507,  -13'd367,  
13'd696,  13'd282,  13'd1027,  13'd213,  -13'd558,  -13'd74,  -13'd168,  13'd179,  -13'd749,  -13'd648,  -13'd794,  -13'd331,  13'd269,  -13'd105,  13'd415,  -13'd129,  
13'd422,  -13'd315,  13'd396,  13'd22,  -13'd495,  13'd272,  -13'd24,  13'd149,  -13'd120,  13'd315,  13'd260,  -13'd14,  -13'd457,  -13'd342,  -13'd246,  -13'd195,  
13'd275,  13'd355,  13'd339,  13'd151,  -13'd247,  -13'd197,  13'd788,  -13'd48,  -13'd247,  -13'd226,  13'd274,  -13'd557,  -13'd763,  13'd760,  13'd566,  13'd694,  
-13'd209,  13'd295,  -13'd189,  -13'd729,  -13'd376,  -13'd48,  13'd114,  -13'd21,  13'd201,  -13'd428,  -13'd385,  -13'd335,  -13'd709,  13'd241,  13'd858,  13'd427,  
13'd527,  -13'd664,  13'd291,  13'd485,  -13'd240,  -13'd193,  -13'd141,  -13'd585,  -13'd642,  13'd437,  -13'd538,  13'd199,  -13'd404,  13'd155,  13'd196,  -13'd30,  
13'd17,  -13'd231,  13'd418,  13'd57,  -13'd343,  13'd524,  13'd70,  13'd171,  13'd377,  -13'd336,  -13'd228,  13'd71,  -13'd278,  13'd146,  -13'd111,  -13'd227,  
-13'd680,  13'd0,  -13'd16,  -13'd269,  -13'd256,  -13'd214,  13'd370,  -13'd483,  -13'd514,  -13'd348,  13'd161,  13'd422,  -13'd302,  -13'd342,  -13'd155,  -13'd906,  
-13'd638,  13'd345,  13'd330,  13'd138,  -13'd352,  13'd382,  13'd381,  -13'd262,  -13'd195,  -13'd432,  -13'd337,  -13'd249,  -13'd69,  13'd615,  13'd516,  13'd229,  
-13'd818,  -13'd473,  13'd453,  13'd25,  -13'd797,  13'd650,  13'd526,  -13'd18,  -13'd389,  13'd107,  13'd542,  13'd312,  13'd44,  13'd4,  13'd248,  -13'd489,  
13'd982,  -13'd1146,  13'd1039,  13'd510,  -13'd500,  13'd831,  -13'd331,  13'd10,  -13'd20,  -13'd26,  13'd1001,  -13'd466,  13'd314,  13'd91,  -13'd251,  13'd348,  
13'd537,  -13'd259,  -13'd792,  13'd233,  -13'd135,  -13'd184,  13'd9,  13'd943,  -13'd332,  13'd132,  -13'd608,  13'd177,  -13'd2,  -13'd566,  -13'd200,  -13'd353,  

-13'd279,  -13'd118,  -13'd84,  -13'd62,  -13'd364,  -13'd235,  -13'd767,  -13'd130,  13'd253,  13'd262,  -13'd96,  13'd73,  13'd107,  13'd578,  13'd216,  -13'd103,  
-13'd506,  -13'd82,  -13'd88,  13'd370,  13'd337,  13'd82,  13'd424,  13'd276,  -13'd57,  -13'd626,  13'd381,  13'd227,  13'd297,  13'd149,  13'd656,  -13'd143,  
-13'd394,  13'd276,  13'd63,  -13'd365,  -13'd540,  13'd31,  13'd283,  -13'd871,  13'd34,  13'd260,  13'd285,  13'd577,  -13'd167,  13'd607,  -13'd115,  -13'd130,  
13'd241,  -13'd520,  -13'd282,  -13'd672,  13'd654,  -13'd139,  13'd45,  13'd399,  13'd384,  -13'd92,  -13'd379,  13'd518,  -13'd111,  -13'd236,  13'd357,  -13'd212,  
-13'd288,  -13'd83,  -13'd275,  -13'd110,  13'd82,  13'd37,  -13'd376,  13'd200,  -13'd550,  13'd401,  -13'd169,  -13'd398,  13'd381,  -13'd497,  13'd1,  13'd335,  
-13'd407,  -13'd213,  -13'd546,  13'd392,  13'd208,  -13'd376,  -13'd201,  -13'd11,  13'd611,  13'd144,  13'd245,  13'd303,  13'd430,  -13'd177,  -13'd247,  -13'd390,  
-13'd590,  -13'd304,  13'd81,  -13'd184,  -13'd19,  -13'd481,  -13'd399,  13'd488,  13'd48,  -13'd417,  13'd38,  -13'd298,  13'd413,  13'd79,  -13'd141,  -13'd187,  
-13'd32,  -13'd346,  -13'd446,  -13'd77,  13'd103,  -13'd296,  -13'd140,  13'd147,  -13'd665,  13'd32,  -13'd455,  -13'd323,  -13'd26,  -13'd606,  -13'd57,  13'd318,  
-13'd359,  -13'd591,  13'd259,  13'd383,  -13'd376,  -13'd133,  -13'd90,  -13'd385,  13'd722,  13'd153,  -13'd137,  -13'd399,  -13'd315,  13'd107,  -13'd13,  13'd0,  
-13'd258,  -13'd300,  -13'd73,  13'd461,  -13'd340,  -13'd209,  13'd649,  -13'd385,  13'd229,  -13'd43,  -13'd123,  -13'd604,  13'd177,  13'd439,  -13'd159,  -13'd89,  
13'd583,  -13'd548,  -13'd736,  13'd213,  -13'd331,  13'd450,  -13'd399,  -13'd500,  13'd529,  -13'd343,  -13'd931,  -13'd448,  -13'd524,  -13'd565,  13'd466,  -13'd229,  
-13'd56,  -13'd854,  13'd222,  13'd362,  13'd537,  -13'd114,  13'd62,  -13'd79,  -13'd460,  13'd567,  13'd364,  -13'd30,  -13'd81,  13'd314,  -13'd49,  -13'd135,  
13'd452,  -13'd283,  -13'd302,  -13'd157,  -13'd227,  13'd36,  -13'd670,  -13'd416,  -13'd383,  -13'd262,  -13'd493,  13'd182,  13'd235,  13'd175,  13'd41,  -13'd97,  
-13'd317,  -13'd606,  13'd155,  -13'd386,  -13'd412,  -13'd756,  -13'd755,  13'd41,  -13'd92,  -13'd333,  13'd605,  -13'd385,  -13'd48,  -13'd367,  -13'd319,  13'd21,  
13'd233,  -13'd160,  -13'd492,  -13'd200,  13'd325,  -13'd544,  13'd397,  13'd23,  -13'd27,  -13'd87,  -13'd156,  -13'd445,  13'd120,  -13'd162,  -13'd150,  13'd42,  
13'd424,  -13'd533,  -13'd507,  -13'd65,  13'd353,  -13'd358,  13'd331,  13'd194,  -13'd22,  13'd571,  -13'd111,  -13'd180,  -13'd284,  -13'd605,  -13'd326,  -13'd140,  
-13'd276,  -13'd149,  -13'd711,  13'd70,  -13'd509,  -13'd300,  -13'd375,  -13'd243,  -13'd179,  -13'd339,  -13'd251,  13'd33,  13'd76,  -13'd438,  -13'd457,  13'd460,  
13'd69,  -13'd232,  13'd241,  -13'd622,  13'd557,  -13'd56,  -13'd848,  -13'd34,  -13'd49,  -13'd799,  -13'd7,  -13'd340,  13'd465,  -13'd374,  -13'd176,  -13'd222,  
13'd46,  13'd355,  13'd493,  -13'd301,  -13'd681,  -13'd526,  -13'd56,  13'd143,  13'd505,  -13'd41,  13'd338,  -13'd260,  13'd301,  13'd605,  -13'd211,  13'd409,  
13'd21,  -13'd662,  13'd328,  13'd268,  -13'd75,  -13'd548,  -13'd273,  13'd725,  -13'd581,  -13'd820,  -13'd484,  13'd129,  -13'd187,  -13'd598,  13'd192,  -13'd94,  
13'd483,  -13'd195,  -13'd515,  -13'd167,  13'd55,  13'd56,  13'd247,  -13'd259,  13'd364,  -13'd18,  13'd44,  13'd67,  13'd191,  -13'd589,  -13'd290,  13'd36,  
13'd239,  13'd275,  -13'd340,  13'd572,  -13'd726,  13'd527,  -13'd133,  -13'd476,  -13'd236,  -13'd193,  -13'd326,  -13'd347,  13'd373,  -13'd81,  13'd286,  13'd317,  
13'd14,  -13'd832,  13'd33,  13'd151,  -13'd241,  -13'd46,  -13'd94,  13'd345,  13'd3,  -13'd312,  13'd535,  -13'd865,  13'd220,  13'd432,  -13'd276,  -13'd262,  
13'd336,  13'd47,  -13'd441,  -13'd201,  13'd416,  -13'd690,  -13'd334,  -13'd275,  13'd392,  -13'd770,  -13'd545,  13'd330,  13'd345,  13'd139,  13'd189,  13'd487,  
-13'd799,  -13'd194,  -13'd749,  13'd23,  -13'd652,  13'd179,  -13'd710,  -13'd192,  13'd436,  -13'd326,  -13'd52,  13'd545,  -13'd91,  -13'd375,  -13'd745,  -13'd185,  

13'd121,  13'd234,  -13'd249,  13'd78,  13'd401,  13'd655,  -13'd243,  -13'd343,  -13'd634,  13'd198,  13'd863,  -13'd420,  13'd742,  -13'd96,  -13'd716,  13'd7,  
-13'd195,  -13'd193,  -13'd832,  13'd909,  -13'd45,  -13'd756,  -13'd1302,  13'd0,  13'd405,  13'd74,  -13'd307,  -13'd220,  13'd347,  -13'd1595,  13'd209,  13'd201,  
-13'd189,  13'd826,  13'd628,  13'd925,  13'd250,  -13'd46,  -13'd500,  -13'd329,  13'd208,  13'd522,  13'd13,  13'd369,  -13'd559,  -13'd823,  13'd815,  13'd105,  
13'd73,  13'd46,  13'd343,  -13'd260,  -13'd102,  13'd85,  13'd255,  -13'd499,  -13'd132,  13'd125,  -13'd159,  13'd693,  13'd451,  13'd1171,  13'd186,  -13'd104,  
-13'd870,  -13'd630,  13'd20,  -13'd88,  13'd73,  -13'd389,  13'd133,  13'd136,  13'd987,  -13'd165,  13'd69,  13'd732,  -13'd821,  -13'd417,  -13'd618,  -13'd501,  
13'd125,  13'd350,  -13'd539,  13'd150,  13'd378,  -13'd386,  -13'd393,  -13'd399,  13'd158,  13'd41,  -13'd49,  -13'd214,  13'd153,  -13'd1194,  13'd324,  13'd366,  
-13'd642,  13'd369,  -13'd837,  -13'd400,  13'd763,  13'd230,  13'd505,  -13'd369,  -13'd50,  13'd561,  -13'd117,  13'd224,  -13'd243,  -13'd1009,  -13'd114,  -13'd391,  
13'd110,  13'd443,  -13'd37,  -13'd51,  13'd402,  13'd48,  -13'd470,  13'd237,  -13'd1026,  -13'd8,  13'd25,  13'd338,  -13'd62,  13'd313,  -13'd687,  13'd1145,  
13'd291,  -13'd26,  13'd140,  -13'd842,  13'd315,  13'd771,  13'd954,  -13'd928,  -13'd744,  -13'd293,  -13'd112,  13'd539,  13'd219,  13'd825,  -13'd565,  13'd743,  
13'd19,  13'd49,  13'd25,  -13'd427,  13'd311,  13'd249,  13'd670,  -13'd159,  -13'd565,  -13'd1155,  13'd168,  -13'd495,  13'd127,  13'd682,  13'd231,  -13'd545,  
-13'd323,  13'd437,  -13'd748,  -13'd94,  13'd529,  13'd303,  -13'd314,  -13'd58,  13'd913,  -13'd275,  13'd384,  13'd267,  -13'd511,  -13'd403,  13'd62,  13'd405,  
-13'd199,  -13'd244,  -13'd495,  13'd261,  13'd879,  13'd210,  -13'd301,  -13'd474,  13'd124,  13'd520,  -13'd698,  -13'd341,  -13'd88,  -13'd199,  13'd298,  13'd163,  
13'd288,  -13'd181,  13'd309,  -13'd84,  -13'd494,  -13'd146,  -13'd620,  13'd285,  13'd168,  -13'd355,  -13'd255,  13'd347,  13'd618,  -13'd168,  13'd793,  -13'd462,  
13'd323,  13'd159,  13'd378,  13'd470,  -13'd200,  -13'd87,  13'd118,  -13'd695,  13'd551,  13'd52,  13'd328,  13'd596,  13'd478,  13'd23,  -13'd270,  13'd148,  
13'd472,  -13'd163,  13'd115,  13'd574,  13'd438,  -13'd256,  13'd373,  13'd116,  13'd77,  13'd271,  -13'd301,  13'd274,  13'd1167,  13'd175,  -13'd630,  13'd114,  
-13'd342,  13'd148,  -13'd848,  -13'd346,  13'd17,  -13'd188,  -13'd118,  -13'd418,  -13'd60,  13'd318,  13'd489,  13'd211,  -13'd125,  -13'd441,  13'd319,  13'd25,  
13'd151,  13'd140,  -13'd22,  -13'd142,  13'd101,  13'd123,  -13'd432,  -13'd734,  13'd1176,  -13'd357,  13'd67,  13'd482,  13'd752,  -13'd639,  -13'd218,  -13'd130,  
-13'd433,  13'd748,  13'd504,  -13'd221,  13'd109,  13'd235,  -13'd271,  13'd280,  13'd84,  13'd567,  -13'd18,  -13'd580,  13'd562,  -13'd975,  -13'd303,  13'd769,  
-13'd345,  -13'd554,  -13'd832,  13'd53,  13'd33,  13'd108,  13'd86,  13'd527,  13'd36,  -13'd93,  13'd819,  13'd218,  13'd516,  -13'd661,  -13'd216,  -13'd548,  
-13'd273,  13'd630,  -13'd814,  13'd234,  13'd429,  -13'd775,  -13'd329,  -13'd150,  13'd307,  13'd1050,  13'd242,  -13'd153,  13'd446,  -13'd149,  13'd492,  -13'd389,  
-13'd24,  -13'd640,  -13'd244,  -13'd375,  -13'd117,  13'd496,  -13'd458,  -13'd312,  13'd499,  -13'd63,  13'd285,  13'd355,  -13'd125,  -13'd222,  13'd877,  -13'd19,  
13'd436,  13'd419,  13'd323,  -13'd20,  13'd93,  -13'd279,  -13'd490,  13'd193,  13'd107,  -13'd424,  13'd180,  13'd289,  13'd191,  13'd165,  -13'd68,  13'd293,  
13'd135,  -13'd233,  -13'd178,  -13'd21,  13'd636,  13'd164,  -13'd405,  -13'd309,  -13'd307,  13'd548,  -13'd300,  13'd682,  -13'd758,  13'd70,  13'd157,  13'd508,  
-13'd131,  13'd525,  13'd312,  13'd84,  13'd538,  13'd742,  13'd295,  13'd303,  -13'd34,  -13'd276,  -13'd335,  13'd262,  -13'd40,  13'd359,  13'd195,  -13'd238,  
-13'd299,  -13'd392,  13'd177,  13'd414,  13'd52,  -13'd331,  13'd467,  -13'd393,  -13'd12,  13'd899,  -13'd380,  13'd158,  13'd386,  13'd31,  -13'd507,  13'd215,  

13'd420,  -13'd326,  13'd484,  -13'd629,  -13'd807,  -13'd377,  -13'd82,  13'd166,  13'd720,  13'd420,  -13'd167,  13'd600,  -13'd80,  -13'd50,  13'd118,  -13'd436,  
13'd419,  -13'd117,  -13'd380,  13'd352,  -13'd501,  -13'd112,  13'd284,  13'd646,  13'd65,  -13'd555,  -13'd339,  13'd355,  -13'd55,  -13'd117,  -13'd372,  -13'd95,  
-13'd685,  -13'd9,  -13'd368,  13'd187,  13'd125,  13'd218,  13'd174,  -13'd54,  -13'd514,  13'd144,  -13'd519,  13'd652,  -13'd7,  13'd216,  -13'd315,  -13'd359,  
-13'd18,  13'd176,  13'd356,  -13'd779,  -13'd39,  -13'd20,  13'd510,  13'd261,  13'd141,  13'd710,  -13'd251,  13'd716,  -13'd387,  -13'd310,  13'd198,  -13'd305,  
13'd647,  13'd53,  13'd943,  13'd187,  -13'd629,  13'd385,  -13'd643,  13'd549,  -13'd303,  13'd541,  13'd315,  13'd320,  -13'd257,  -13'd340,  13'd490,  13'd750,  
13'd192,  -13'd289,  -13'd28,  -13'd6,  13'd360,  -13'd24,  -13'd505,  13'd864,  13'd932,  13'd761,  -13'd514,  13'd351,  13'd295,  13'd139,  13'd659,  -13'd507,  
-13'd406,  -13'd450,  -13'd38,  13'd408,  -13'd73,  13'd108,  13'd473,  13'd465,  13'd651,  -13'd45,  13'd181,  13'd31,  13'd238,  13'd41,  13'd45,  -13'd48,  
-13'd99,  -13'd373,  13'd186,  13'd114,  -13'd479,  13'd346,  -13'd321,  13'd59,  13'd128,  13'd273,  -13'd127,  13'd339,  13'd654,  -13'd403,  13'd57,  13'd239,  
-13'd421,  13'd506,  13'd327,  -13'd146,  -13'd169,  -13'd350,  13'd93,  13'd290,  13'd124,  -13'd483,  -13'd272,  13'd43,  13'd336,  -13'd176,  13'd72,  13'd364,  
13'd912,  -13'd15,  13'd493,  -13'd2,  13'd268,  -13'd745,  -13'd505,  13'd382,  -13'd311,  13'd110,  13'd343,  13'd186,  13'd945,  13'd31,  -13'd120,  13'd1007,  
13'd232,  13'd625,  13'd160,  13'd181,  13'd1162,  13'd412,  -13'd286,  13'd790,  -13'd122,  -13'd802,  -13'd288,  -13'd87,  13'd836,  13'd492,  -13'd311,  13'd244,  
-13'd61,  13'd236,  13'd694,  13'd807,  13'd241,  -13'd138,  13'd795,  13'd97,  13'd333,  -13'd970,  13'd256,  -13'd385,  13'd29,  13'd124,  -13'd452,  13'd270,  
-13'd122,  13'd407,  -13'd149,  -13'd132,  -13'd98,  13'd466,  13'd109,  -13'd24,  13'd274,  -13'd820,  13'd388,  13'd226,  -13'd4,  -13'd1083,  13'd198,  -13'd180,  
13'd379,  -13'd83,  -13'd579,  13'd168,  -13'd405,  -13'd815,  -13'd523,  13'd108,  -13'd855,  -13'd738,  13'd0,  13'd348,  13'd471,  13'd941,  13'd329,  -13'd538,  
13'd954,  -13'd72,  -13'd57,  13'd568,  -13'd96,  13'd351,  13'd399,  -13'd351,  -13'd507,  -13'd536,  13'd3,  -13'd326,  13'd1014,  -13'd439,  -13'd339,  13'd529,  
13'd104,  13'd367,  -13'd473,  -13'd376,  -13'd120,  13'd541,  -13'd286,  -13'd181,  -13'd638,  -13'd491,  -13'd631,  13'd979,  -13'd36,  -13'd84,  -13'd349,  -13'd383,  
-13'd104,  -13'd150,  -13'd261,  -13'd198,  13'd380,  -13'd479,  -13'd414,  -13'd68,  13'd70,  13'd361,  -13'd834,  -13'd23,  -13'd101,  13'd489,  13'd214,  13'd512,  
-13'd755,  13'd650,  -13'd358,  -13'd109,  13'd103,  -13'd52,  13'd84,  -13'd766,  -13'd280,  -13'd329,  13'd343,  13'd20,  -13'd290,  -13'd294,  -13'd58,  13'd244,  
-13'd48,  -13'd278,  -13'd393,  -13'd169,  13'd47,  13'd576,  -13'd461,  13'd70,  -13'd257,  13'd223,  13'd343,  13'd87,  13'd472,  13'd34,  13'd62,  13'd391,  
-13'd393,  -13'd118,  13'd1222,  -13'd585,  13'd219,  -13'd193,  13'd17,  13'd256,  -13'd247,  13'd44,  13'd320,  13'd165,  13'd442,  13'd285,  -13'd457,  -13'd386,  
13'd386,  13'd851,  13'd588,  -13'd147,  13'd62,  -13'd124,  -13'd1251,  -13'd5,  -13'd830,  13'd428,  -13'd230,  13'd508,  13'd430,  13'd400,  13'd275,  -13'd738,  
13'd10,  -13'd439,  -13'd481,  -13'd97,  -13'd96,  -13'd686,  -13'd962,  -13'd43,  -13'd521,  13'd150,  -13'd565,  -13'd4,  -13'd277,  13'd572,  13'd351,  13'd215,  
-13'd284,  13'd59,  -13'd23,  -13'd216,  13'd135,  -13'd83,  13'd185,  13'd120,  -13'd734,  -13'd1007,  -13'd263,  -13'd70,  -13'd290,  -13'd295,  -13'd241,  -13'd387,  
13'd913,  -13'd371,  -13'd283,  -13'd25,  13'd5,  13'd171,  -13'd574,  -13'd365,  -13'd46,  -13'd262,  -13'd139,  13'd674,  13'd50,  13'd857,  13'd228,  -13'd56,  
13'd248,  -13'd74,  13'd512,  13'd584,  13'd299,  -13'd13,  13'd465,  -13'd412,  -13'd223,  -13'd1225,  -13'd710,  13'd195,  13'd336,  13'd209,  -13'd388,  -13'd250,  

-13'd505,  13'd32,  13'd221,  13'd190,  13'd345,  13'd350,  -13'd1294,  13'd30,  -13'd68,  -13'd104,  -13'd311,  13'd489,  -13'd109,  13'd70,  13'd139,  -13'd159,  
13'd325,  -13'd184,  -13'd22,  -13'd546,  13'd39,  -13'd2,  13'd346,  -13'd110,  13'd284,  -13'd373,  -13'd134,  -13'd114,  13'd681,  -13'd767,  13'd601,  -13'd139,  
-13'd329,  13'd457,  13'd228,  13'd206,  -13'd331,  -13'd355,  -13'd118,  13'd173,  13'd283,  -13'd831,  -13'd693,  -13'd146,  13'd388,  13'd221,  13'd192,  13'd187,  
13'd67,  13'd1078,  13'd81,  -13'd482,  13'd415,  13'd112,  -13'd814,  -13'd47,  13'd679,  13'd432,  -13'd856,  -13'd362,  13'd168,  -13'd271,  13'd706,  13'd571,  
13'd679,  -13'd280,  13'd436,  13'd429,  -13'd232,  13'd27,  -13'd819,  13'd351,  13'd246,  13'd512,  -13'd540,  13'd89,  -13'd397,  -13'd450,  -13'd69,  -13'd1342,  
-13'd307,  13'd736,  13'd188,  -13'd99,  13'd304,  13'd116,  13'd652,  -13'd410,  13'd25,  -13'd362,  13'd116,  -13'd146,  13'd386,  13'd496,  13'd147,  13'd353,  
13'd193,  -13'd165,  -13'd469,  13'd438,  13'd198,  13'd108,  13'd957,  13'd169,  13'd28,  -13'd455,  13'd648,  13'd96,  13'd34,  -13'd884,  -13'd451,  13'd22,  
-13'd697,  13'd1188,  -13'd478,  -13'd29,  13'd415,  13'd43,  13'd322,  13'd223,  -13'd86,  -13'd159,  -13'd337,  13'd215,  13'd83,  13'd138,  -13'd835,  -13'd321,  
-13'd567,  13'd1584,  -13'd94,  13'd429,  13'd520,  -13'd617,  -13'd256,  -13'd75,  13'd395,  -13'd147,  13'd9,  13'd658,  13'd133,  -13'd241,  13'd591,  13'd244,  
13'd895,  13'd906,  13'd818,  -13'd381,  13'd558,  13'd320,  13'd65,  -13'd771,  -13'd338,  -13'd152,  13'd129,  13'd307,  13'd272,  -13'd250,  13'd327,  13'd251,  
13'd580,  13'd482,  13'd407,  13'd382,  -13'd229,  13'd374,  13'd141,  13'd141,  -13'd575,  -13'd548,  -13'd477,  13'd724,  13'd428,  13'd198,  -13'd134,  13'd431,  
-13'd194,  -13'd32,  -13'd224,  13'd74,  13'd344,  -13'd267,  13'd401,  13'd213,  13'd925,  -13'd1025,  -13'd163,  -13'd271,  -13'd536,  -13'd350,  -13'd181,  13'd120,  
-13'd457,  13'd218,  13'd313,  13'd410,  13'd810,  -13'd848,  13'd78,  13'd316,  -13'd314,  13'd114,  -13'd44,  13'd214,  -13'd649,  13'd186,  -13'd103,  -13'd22,  
13'd512,  -13'd20,  -13'd182,  13'd527,  -13'd771,  13'd517,  -13'd173,  13'd280,  -13'd309,  -13'd442,  13'd185,  13'd324,  -13'd208,  13'd639,  13'd399,  13'd388,  
13'd1174,  13'd583,  13'd381,  -13'd36,  -13'd1091,  13'd103,  13'd789,  13'd339,  13'd258,  -13'd112,  -13'd161,  13'd406,  -13'd225,  -13'd147,  13'd790,  -13'd566,  
-13'd105,  -13'd193,  -13'd41,  13'd108,  -13'd315,  -13'd198,  13'd630,  13'd15,  -13'd570,  -13'd539,  -13'd112,  -13'd433,  -13'd623,  -13'd223,  13'd48,  -13'd410,  
13'd451,  13'd10,  -13'd782,  13'd690,  13'd117,  13'd195,  13'd392,  -13'd338,  13'd362,  -13'd211,  -13'd739,  -13'd58,  -13'd420,  -13'd562,  13'd714,  13'd73,  
13'd190,  13'd319,  -13'd358,  13'd60,  -13'd137,  13'd426,  13'd644,  -13'd181,  13'd681,  13'd588,  13'd44,  -13'd373,  -13'd159,  -13'd194,  -13'd106,  -13'd824,  
13'd681,  13'd653,  13'd766,  13'd218,  -13'd80,  13'd696,  13'd13,  13'd341,  -13'd155,  13'd359,  13'd170,  -13'd147,  13'd386,  -13'd276,  13'd229,  -13'd58,  
13'd188,  -13'd15,  -13'd186,  13'd221,  13'd89,  13'd197,  -13'd29,  13'd130,  13'd95,  -13'd293,  13'd162,  -13'd430,  13'd662,  -13'd497,  13'd156,  13'd739,  
13'd176,  13'd210,  13'd443,  -13'd200,  -13'd474,  -13'd766,  -13'd789,  -13'd348,  -13'd1008,  13'd532,  -13'd1362,  13'd119,  -13'd298,  13'd0,  -13'd327,  -13'd711,  
13'd478,  13'd379,  13'd837,  13'd79,  -13'd232,  13'd968,  -13'd22,  -13'd205,  -13'd151,  13'd475,  -13'd310,  -13'd186,  13'd40,  13'd799,  13'd196,  13'd155,  
-13'd383,  -13'd200,  -13'd106,  13'd352,  -13'd110,  13'd85,  -13'd506,  13'd184,  13'd85,  -13'd39,  13'd101,  -13'd283,  13'd480,  -13'd322,  13'd3,  -13'd674,  
-13'd805,  -13'd519,  -13'd468,  -13'd201,  13'd968,  13'd3,  13'd464,  13'd379,  -13'd1177,  13'd449,  -13'd679,  -13'd91,  -13'd226,  -13'd348,  13'd663,  13'd291,  
-13'd874,  -13'd205,  -13'd1232,  13'd425,  13'd382,  13'd33,  -13'd193,  13'd196,  -13'd663,  -13'd157,  -13'd106,  -13'd517,  -13'd546,  -13'd337,  -13'd353,  13'd37,  

-13'd478,  13'd1096,  -13'd423,  -13'd33,  13'd619,  13'd653,  -13'd362,  13'd341,  -13'd867,  -13'd310,  -13'd200,  -13'd81,  13'd455,  -13'd252,  13'd146,  13'd410,  
13'd173,  13'd927,  -13'd464,  -13'd4,  13'd672,  13'd1052,  -13'd916,  -13'd546,  -13'd257,  13'd339,  -13'd207,  13'd56,  13'd34,  13'd210,  13'd636,  13'd977,  
-13'd28,  13'd65,  13'd369,  -13'd529,  13'd413,  -13'd297,  13'd1044,  13'd25,  -13'd162,  -13'd420,  13'd16,  13'd422,  13'd230,  13'd921,  -13'd480,  -13'd100,  
-13'd509,  -13'd432,  13'd498,  -13'd56,  -13'd867,  -13'd213,  -13'd123,  -13'd390,  13'd629,  13'd45,  13'd475,  13'd22,  -13'd559,  13'd859,  -13'd449,  13'd293,  
-13'd1145,  -13'd1219,  13'd413,  -13'd61,  -13'd666,  -13'd715,  13'd21,  -13'd517,  -13'd10,  -13'd388,  -13'd196,  -13'd659,  -13'd915,  -13'd388,  13'd202,  -13'd50,  
-13'd17,  -13'd254,  13'd214,  13'd21,  -13'd228,  -13'd227,  -13'd569,  13'd564,  -13'd553,  -13'd32,  13'd345,  13'd318,  13'd488,  -13'd481,  -13'd623,  13'd874,  
13'd627,  13'd1310,  -13'd780,  -13'd56,  13'd142,  13'd180,  -13'd280,  13'd422,  13'd295,  -13'd479,  -13'd634,  13'd181,  13'd356,  13'd448,  13'd323,  13'd464,  
13'd221,  13'd68,  -13'd216,  -13'd90,  -13'd457,  -13'd215,  13'd877,  -13'd28,  -13'd231,  -13'd559,  13'd366,  13'd236,  13'd299,  13'd419,  -13'd16,  13'd205,  
13'd471,  13'd83,  13'd903,  -13'd789,  13'd384,  -13'd109,  13'd872,  13'd228,  13'd278,  13'd199,  13'd109,  13'd349,  -13'd959,  13'd843,  -13'd680,  13'd317,  
13'd63,  -13'd27,  13'd797,  13'd58,  -13'd231,  13'd33,  13'd499,  13'd563,  -13'd237,  -13'd288,  -13'd447,  13'd517,  13'd217,  -13'd967,  -13'd669,  -13'd811,  
-13'd463,  13'd325,  -13'd365,  13'd186,  -13'd141,  -13'd505,  -13'd769,  -13'd218,  -13'd289,  -13'd338,  13'd839,  -13'd381,  -13'd460,  13'd51,  13'd51,  13'd84,  
13'd909,  13'd103,  -13'd227,  -13'd154,  -13'd568,  13'd364,  -13'd846,  -13'd5,  -13'd131,  -13'd240,  -13'd718,  13'd740,  -13'd318,  13'd179,  -13'd95,  -13'd492,  
-13'd58,  13'd23,  13'd521,  -13'd494,  -13'd171,  13'd355,  13'd400,  13'd874,  13'd477,  -13'd708,  13'd21,  -13'd391,  -13'd184,  -13'd59,  13'd121,  13'd446,  
-13'd332,  13'd533,  -13'd72,  13'd738,  13'd481,  13'd79,  13'd270,  13'd72,  13'd195,  13'd318,  -13'd330,  -13'd569,  13'd90,  -13'd9,  -13'd403,  -13'd402,  
-13'd38,  -13'd695,  13'd382,  13'd494,  -13'd155,  -13'd27,  -13'd917,  -13'd69,  13'd631,  13'd357,  13'd242,  13'd596,  -13'd219,  -13'd375,  13'd321,  13'd621,  
13'd0,  -13'd30,  13'd516,  13'd526,  -13'd671,  13'd60,  13'd271,  13'd560,  13'd519,  -13'd350,  13'd492,  -13'd611,  -13'd45,  13'd269,  -13'd244,  -13'd458,  
13'd548,  -13'd576,  13'd393,  -13'd138,  13'd482,  13'd78,  13'd985,  -13'd106,  -13'd256,  -13'd760,  13'd641,  -13'd54,  -13'd660,  -13'd382,  13'd224,  13'd409,  
13'd7,  13'd59,  -13'd97,  -13'd506,  -13'd108,  13'd60,  -13'd263,  13'd179,  13'd162,  -13'd367,  -13'd181,  -13'd478,  -13'd148,  -13'd81,  -13'd711,  13'd102,  
13'd53,  -13'd313,  -13'd982,  -13'd3,  -13'd35,  -13'd288,  -13'd1139,  13'd158,  13'd432,  13'd344,  -13'd726,  13'd319,  -13'd96,  13'd778,  13'd461,  13'd885,  
13'd492,  13'd293,  13'd603,  13'd317,  13'd393,  13'd834,  13'd400,  -13'd190,  13'd464,  13'd1032,  13'd396,  13'd336,  13'd75,  -13'd795,  13'd265,  13'd213,  
13'd361,  -13'd82,  13'd65,  13'd458,  -13'd215,  13'd750,  13'd619,  13'd214,  13'd516,  13'd539,  13'd471,  -13'd79,  13'd264,  -13'd163,  13'd90,  -13'd239,  
13'd366,  -13'd89,  13'd14,  13'd104,  -13'd157,  -13'd551,  -13'd252,  -13'd77,  -13'd36,  -13'd755,  -13'd135,  -13'd764,  13'd390,  13'd173,  -13'd759,  -13'd196,  
-13'd667,  -13'd258,  -13'd343,  -13'd311,  13'd685,  -13'd515,  -13'd465,  -13'd14,  -13'd740,  13'd850,  -13'd164,  13'd461,  13'd563,  -13'd393,  13'd129,  -13'd132,  
13'd124,  13'd302,  -13'd141,  -13'd834,  -13'd316,  13'd99,  -13'd1182,  -13'd399,  13'd1061,  13'd931,  -13'd415,  13'd320,  -13'd62,  -13'd466,  -13'd460,  13'd22,  
13'd473,  -13'd14,  13'd30,  -13'd212,  -13'd5,  13'd656,  -13'd65,  -13'd10,  13'd229,  13'd182,  13'd53,  13'd481,  13'd976,  -13'd120,  13'd521,  -13'd85,  

-13'd923,  -13'd1303,  -13'd655,  -13'd880,  13'd464,  -13'd557,  13'd598,  -13'd510,  -13'd573,  13'd544,  -13'd930,  -13'd105,  -13'd235,  -13'd90,  -13'd1086,  -13'd1110,  
13'd193,  13'd516,  -13'd72,  -13'd651,  -13'd704,  -13'd512,  -13'd223,  -13'd9,  -13'd1022,  -13'd342,  -13'd452,  -13'd296,  -13'd275,  13'd981,  -13'd631,  -13'd519,  
13'd1229,  -13'd95,  13'd1067,  13'd527,  -13'd486,  13'd357,  13'd539,  -13'd204,  -13'd242,  -13'd822,  -13'd8,  13'd12,  13'd63,  13'd888,  -13'd530,  -13'd522,  
13'd342,  -13'd5,  -13'd150,  13'd284,  -13'd603,  -13'd373,  13'd215,  13'd54,  13'd232,  -13'd94,  13'd700,  13'd447,  -13'd363,  -13'd702,  -13'd28,  -13'd42,  
13'd222,  13'd156,  13'd104,  13'd182,  -13'd265,  -13'd287,  -13'd66,  13'd307,  -13'd611,  13'd400,  -13'd103,  13'd299,  13'd144,  -13'd268,  13'd277,  13'd693,  
-13'd925,  -13'd64,  -13'd1349,  -13'd170,  13'd73,  -13'd272,  -13'd438,  13'd23,  13'd476,  13'd125,  13'd23,  -13'd138,  -13'd25,  -13'd678,  -13'd69,  -13'd112,  
13'd335,  13'd294,  13'd391,  13'd397,  13'd404,  -13'd211,  -13'd866,  -13'd735,  -13'd730,  -13'd623,  13'd659,  13'd461,  -13'd81,  13'd1043,  -13'd288,  -13'd253,  
13'd689,  -13'd11,  13'd608,  -13'd76,  -13'd730,  -13'd103,  -13'd397,  13'd521,  13'd422,  13'd554,  -13'd447,  13'd174,  -13'd671,  13'd502,  -13'd551,  -13'd155,  
-13'd70,  13'd425,  13'd42,  -13'd356,  13'd233,  13'd227,  13'd288,  13'd115,  -13'd321,  13'd258,  13'd546,  -13'd174,  13'd239,  13'd696,  13'd515,  -13'd24,  
-13'd6,  -13'd832,  -13'd1111,  13'd275,  -13'd216,  -13'd942,  13'd239,  -13'd129,  13'd667,  -13'd645,  -13'd37,  -13'd75,  -13'd1242,  13'd228,  13'd138,  13'd72,  
-13'd195,  13'd51,  -13'd761,  13'd500,  13'd243,  -13'd520,  -13'd1422,  13'd169,  13'd388,  -13'd108,  13'd481,  -13'd158,  -13'd275,  -13'd954,  13'd483,  13'd30,  
-13'd62,  -13'd383,  -13'd24,  -13'd275,  -13'd795,  -13'd1234,  -13'd128,  -13'd1112,  -13'd392,  13'd381,  -13'd299,  -13'd526,  -13'd70,  13'd898,  -13'd326,  -13'd197,  
13'd529,  -13'd11,  13'd432,  -13'd247,  -13'd217,  -13'd489,  13'd410,  13'd615,  -13'd80,  -13'd106,  -13'd579,  13'd193,  13'd361,  13'd620,  -13'd241,  -13'd18,  
-13'd64,  13'd587,  13'd1112,  -13'd401,  -13'd674,  13'd384,  13'd952,  -13'd287,  13'd552,  -13'd750,  -13'd12,  -13'd4,  -13'd557,  13'd182,  -13'd85,  13'd103,  
13'd785,  13'd614,  -13'd599,  13'd223,  -13'd445,  -13'd893,  13'd328,  13'd696,  -13'd62,  -13'd1388,  13'd539,  -13'd315,  -13'd406,  -13'd674,  13'd481,  -13'd1235,  
-13'd46,  13'd223,  -13'd162,  -13'd129,  13'd694,  13'd143,  -13'd129,  13'd70,  -13'd343,  13'd394,  13'd40,  -13'd1505,  -13'd644,  -13'd420,  -13'd254,  -13'd451,  
-13'd38,  -13'd1183,  -13'd59,  -13'd471,  13'd382,  -13'd619,  13'd559,  -13'd536,  -13'd1720,  13'd523,  13'd162,  13'd83,  13'd555,  13'd60,  13'd606,  -13'd374,  
-13'd12,  -13'd666,  13'd714,  -13'd445,  -13'd1295,  -13'd451,  13'd417,  -13'd547,  13'd326,  -13'd388,  -13'd1334,  -13'd314,  -13'd260,  13'd764,  -13'd109,  -13'd1452,  
13'd104,  13'd104,  13'd1172,  13'd606,  -13'd1255,  -13'd709,  -13'd301,  13'd44,  -13'd50,  13'd624,  -13'd162,  13'd18,  -13'd764,  -13'd384,  13'd244,  -13'd1602,  
13'd159,  13'd323,  -13'd91,  13'd76,  -13'd1599,  -13'd975,  -13'd167,  -13'd48,  -13'd897,  13'd599,  -13'd975,  13'd522,  -13'd129,  -13'd128,  -13'd573,  -13'd983,  
13'd109,  13'd4,  -13'd419,  13'd747,  -13'd331,  -13'd50,  13'd202,  13'd596,  13'd142,  -13'd112,  -13'd375,  -13'd478,  -13'd214,  -13'd522,  13'd10,  13'd386,  
13'd817,  13'd17,  13'd344,  13'd527,  -13'd1586,  13'd580,  -13'd338,  -13'd40,  13'd763,  13'd950,  -13'd469,  -13'd110,  -13'd285,  -13'd229,  13'd1,  13'd223,  
13'd77,  -13'd410,  13'd193,  13'd245,  13'd397,  -13'd133,  13'd492,  -13'd83,  13'd718,  13'd1299,  13'd208,  -13'd24,  -13'd298,  -13'd487,  13'd311,  13'd367,  
-13'd572,  -13'd687,  13'd409,  13'd479,  13'd103,  -13'd834,  -13'd523,  13'd408,  13'd448,  13'd79,  13'd407,  -13'd173,  -13'd67,  13'd227,  13'd314,  13'd903,  
-13'd171,  -13'd562,  -13'd95,  13'd252,  -13'd26,  -13'd920,  13'd109,  13'd89,  -13'd941,  13'd535,  13'd190,  13'd738,  13'd221,  13'd81,  13'd180,  13'd745,  

13'd293,  -13'd166,  -13'd371,  -13'd11,  13'd877,  -13'd579,  13'd522,  -13'd281,  -13'd109,  13'd560,  13'd165,  -13'd50,  -13'd653,  -13'd579,  -13'd280,  13'd425,  
-13'd280,  -13'd72,  -13'd888,  -13'd594,  13'd385,  13'd198,  13'd682,  13'd196,  13'd45,  -13'd219,  -13'd1131,  -13'd95,  13'd692,  13'd171,  -13'd72,  -13'd78,  
-13'd18,  -13'd29,  -13'd315,  -13'd697,  -13'd172,  -13'd19,  -13'd150,  13'd0,  -13'd377,  -13'd662,  -13'd630,  13'd554,  13'd72,  13'd367,  13'd306,  13'd317,  
13'd315,  13'd344,  -13'd621,  -13'd346,  -13'd3,  -13'd14,  13'd518,  -13'd309,  13'd642,  -13'd225,  -13'd38,  13'd136,  13'd254,  13'd1505,  13'd377,  13'd483,  
-13'd195,  -13'd116,  13'd58,  -13'd203,  13'd135,  13'd241,  13'd109,  13'd352,  -13'd102,  -13'd8,  13'd26,  -13'd369,  -13'd483,  13'd251,  13'd865,  13'd261,  
13'd28,  13'd824,  -13'd307,  -13'd474,  -13'd457,  -13'd251,  13'd693,  -13'd764,  -13'd306,  13'd480,  13'd509,  13'd156,  13'd9,  -13'd1033,  -13'd8,  -13'd188,  
13'd473,  13'd483,  -13'd236,  -13'd236,  13'd85,  -13'd155,  -13'd235,  -13'd510,  13'd465,  13'd698,  -13'd146,  -13'd385,  -13'd316,  -13'd436,  -13'd40,  13'd114,  
-13'd86,  13'd621,  13'd46,  -13'd553,  13'd260,  13'd683,  -13'd247,  13'd75,  13'd155,  -13'd146,  13'd239,  -13'd82,  -13'd29,  -13'd42,  -13'd268,  -13'd134,  
13'd445,  13'd1,  13'd669,  13'd363,  13'd274,  13'd239,  13'd495,  13'd51,  -13'd342,  -13'd661,  13'd60,  13'd389,  -13'd163,  13'd156,  -13'd244,  -13'd494,  
13'd20,  13'd450,  13'd631,  13'd608,  -13'd235,  13'd772,  -13'd241,  13'd5,  13'd424,  -13'd289,  13'd151,  -13'd128,  -13'd514,  13'd539,  13'd749,  -13'd731,  
13'd6,  13'd351,  -13'd447,  13'd54,  -13'd685,  13'd235,  13'd397,  -13'd134,  -13'd90,  13'd191,  -13'd594,  13'd978,  13'd241,  -13'd68,  13'd306,  13'd31,  
-13'd78,  -13'd44,  -13'd509,  -13'd229,  -13'd76,  -13'd399,  -13'd144,  13'd47,  13'd1081,  13'd112,  -13'd791,  13'd112,  -13'd612,  -13'd7,  -13'd41,  -13'd465,  
13'd206,  13'd383,  -13'd773,  13'd622,  13'd495,  -13'd552,  13'd279,  13'd48,  13'd146,  13'd27,  -13'd100,  13'd211,  -13'd269,  -13'd60,  -13'd291,  13'd400,  
13'd694,  -13'd61,  13'd311,  13'd180,  -13'd555,  13'd327,  13'd42,  13'd440,  13'd289,  13'd451,  -13'd65,  -13'd79,  -13'd222,  13'd253,  13'd721,  13'd154,  
13'd456,  13'd223,  -13'd118,  13'd293,  -13'd98,  13'd617,  13'd288,  13'd436,  -13'd202,  -13'd223,  -13'd219,  13'd47,  13'd669,  13'd98,  13'd218,  13'd322,  
13'd462,  13'd426,  13'd569,  13'd810,  13'd217,  13'd115,  13'd466,  13'd493,  -13'd346,  13'd320,  13'd100,  -13'd356,  13'd331,  13'd529,  13'd608,  -13'd96,  
13'd578,  -13'd211,  13'd617,  13'd161,  -13'd463,  -13'd214,  -13'd127,  13'd115,  -13'd3,  -13'd691,  -13'd174,  -13'd340,  -13'd379,  13'd134,  13'd457,  -13'd575,  
13'd606,  13'd319,  -13'd1089,  13'd315,  13'd406,  13'd112,  -13'd561,  13'd566,  -13'd950,  -13'd129,  13'd426,  -13'd170,  13'd688,  -13'd161,  -13'd1,  13'd447,  
13'd157,  -13'd573,  13'd87,  -13'd25,  13'd628,  13'd212,  -13'd580,  13'd634,  -13'd581,  13'd57,  -13'd580,  -13'd325,  13'd171,  13'd633,  -13'd227,  13'd905,  
13'd228,  13'd284,  -13'd27,  13'd831,  13'd176,  13'd483,  13'd464,  13'd154,  13'd212,  13'd413,  13'd252,  13'd94,  13'd560,  13'd458,  -13'd0,  -13'd249,  
13'd366,  -13'd104,  13'd331,  13'd954,  13'd1228,  13'd630,  -13'd703,  13'd679,  -13'd745,  13'd209,  13'd48,  13'd82,  13'd761,  13'd125,  13'd810,  13'd64,  
-13'd834,  13'd95,  13'd304,  13'd772,  13'd307,  -13'd59,  -13'd282,  13'd342,  -13'd26,  -13'd125,  -13'd206,  -13'd167,  -13'd261,  13'd755,  13'd397,  -13'd180,  
-13'd474,  13'd626,  -13'd552,  -13'd557,  -13'd313,  -13'd56,  -13'd693,  13'd278,  -13'd1133,  -13'd347,  13'd605,  -13'd24,  -13'd158,  -13'd1067,  -13'd627,  -13'd193,  
13'd244,  -13'd116,  13'd261,  13'd578,  -13'd242,  13'd513,  13'd153,  13'd714,  13'd179,  13'd211,  -13'd309,  13'd443,  -13'd174,  -13'd464,  -13'd727,  -13'd478,  
13'd129,  13'd4,  13'd221,  13'd255,  -13'd391,  13'd404,  13'd344,  13'd147,  13'd790,  13'd29,  13'd69,  13'd84,  13'd619,  -13'd487,  -13'd165,  -13'd103,  

13'd78,  13'd406,  -13'd345,  -13'd777,  13'd62,  -13'd540,  13'd485,  -13'd968,  -13'd725,  -13'd503,  -13'd390,  13'd587,  -13'd216,  13'd144,  -13'd67,  -13'd699,  
13'd316,  -13'd229,  -13'd128,  -13'd350,  -13'd48,  -13'd9,  13'd49,  -13'd461,  -13'd762,  13'd11,  -13'd157,  13'd67,  -13'd377,  13'd273,  13'd225,  13'd602,  
13'd449,  13'd906,  -13'd444,  -13'd210,  13'd381,  -13'd202,  13'd460,  -13'd560,  -13'd127,  13'd484,  13'd314,  13'd420,  -13'd725,  13'd134,  -13'd22,  13'd201,  
13'd700,  -13'd444,  13'd456,  13'd291,  -13'd439,  -13'd353,  13'd347,  -13'd1027,  -13'd248,  13'd646,  13'd295,  -13'd151,  -13'd97,  -13'd94,  13'd422,  13'd246,  
-13'd589,  -13'd1338,  -13'd503,  -13'd667,  -13'd93,  13'd56,  13'd372,  13'd126,  -13'd564,  -13'd685,  -13'd286,  13'd306,  13'd155,  -13'd665,  -13'd563,  13'd437,  
-13'd24,  -13'd210,  13'd260,  -13'd858,  -13'd746,  -13'd252,  13'd182,  -13'd669,  13'd516,  -13'd377,  13'd804,  13'd27,  -13'd922,  13'd149,  -13'd376,  13'd194,  
-13'd134,  13'd484,  -13'd88,  -13'd114,  13'd271,  13'd468,  13'd49,  -13'd418,  -13'd666,  -13'd109,  -13'd529,  13'd118,  -13'd11,  13'd115,  -13'd661,  -13'd738,  
13'd216,  -13'd36,  -13'd365,  13'd247,  -13'd489,  13'd78,  13'd395,  -13'd833,  -13'd200,  -13'd9,  -13'd381,  13'd423,  -13'd430,  -13'd56,  13'd12,  13'd695,  
13'd450,  13'd653,  13'd263,  -13'd1036,  -13'd405,  13'd171,  13'd826,  13'd318,  -13'd281,  13'd892,  13'd28,  13'd166,  13'd219,  13'd799,  -13'd296,  13'd129,  
13'd364,  13'd593,  13'd1056,  -13'd583,  -13'd484,  -13'd648,  13'd176,  -13'd432,  13'd595,  -13'd633,  -13'd130,  -13'd576,  -13'd752,  13'd33,  -13'd543,  13'd310,  
-13'd769,  -13'd529,  13'd726,  13'd407,  -13'd45,  -13'd50,  -13'd205,  13'd294,  13'd380,  13'd455,  -13'd705,  -13'd362,  -13'd517,  -13'd218,  13'd301,  -13'd314,  
13'd41,  13'd219,  -13'd207,  -13'd10,  -13'd650,  13'd155,  13'd466,  13'd258,  -13'd147,  -13'd128,  13'd129,  -13'd392,  13'd241,  -13'd16,  -13'd233,  13'd19,  
13'd741,  13'd181,  13'd1151,  -13'd80,  -13'd753,  13'd730,  13'd562,  13'd317,  -13'd342,  -13'd92,  13'd181,  13'd359,  13'd244,  13'd949,  13'd227,  13'd611,  
13'd595,  13'd774,  13'd892,  -13'd101,  -13'd687,  -13'd321,  13'd827,  13'd1011,  13'd421,  13'd223,  13'd462,  13'd570,  -13'd171,  13'd772,  13'd216,  -13'd620,  
13'd229,  13'd234,  -13'd399,  -13'd310,  13'd83,  -13'd549,  13'd274,  -13'd39,  -13'd485,  -13'd740,  -13'd443,  -13'd288,  13'd255,  13'd258,  -13'd678,  -13'd342,  
13'd484,  -13'd700,  -13'd316,  -13'd538,  -13'd779,  13'd377,  13'd579,  -13'd201,  13'd754,  -13'd45,  13'd620,  -13'd61,  -13'd158,  13'd267,  -13'd181,  -13'd327,  
13'd119,  13'd334,  13'd140,  13'd285,  -13'd192,  -13'd211,  13'd686,  13'd447,  -13'd458,  -13'd409,  13'd1052,  -13'd1,  13'd478,  13'd894,  13'd164,  13'd15,  
-13'd707,  13'd411,  13'd925,  -13'd174,  -13'd398,  13'd198,  13'd805,  13'd228,  13'd317,  13'd352,  -13'd607,  -13'd600,  13'd365,  13'd1250,  -13'd296,  -13'd63,  
-13'd129,  -13'd519,  13'd194,  13'd80,  13'd45,  -13'd927,  -13'd232,  -13'd10,  -13'd888,  -13'd810,  -13'd816,  -13'd32,  -13'd314,  13'd281,  -13'd511,  -13'd346,  
13'd79,  13'd14,  13'd597,  13'd557,  -13'd1201,  -13'd861,  -13'd767,  -13'd425,  -13'd116,  -13'd186,  -13'd491,  -13'd328,  -13'd70,  13'd797,  -13'd164,  -13'd837,  
-13'd622,  13'd455,  -13'd457,  -13'd660,  13'd319,  -13'd67,  13'd1133,  13'd514,  -13'd299,  13'd402,  13'd145,  13'd610,  -13'd275,  -13'd1095,  -13'd254,  13'd209,  
-13'd329,  13'd140,  -13'd245,  13'd226,  13'd622,  -13'd566,  13'd515,  -13'd81,  13'd651,  13'd413,  13'd347,  -13'd778,  -13'd396,  13'd579,  -13'd393,  -13'd655,  
-13'd134,  -13'd153,  13'd633,  13'd11,  13'd451,  -13'd61,  13'd666,  13'd543,  13'd786,  13'd769,  -13'd44,  -13'd1220,  -13'd314,  13'd669,  13'd343,  -13'd525,  
-13'd1025,  -13'd213,  -13'd380,  13'd127,  13'd620,  -13'd368,  -13'd482,  -13'd629,  13'd270,  13'd592,  13'd212,  -13'd292,  13'd126,  13'd401,  13'd94,  -13'd463,  
13'd81,  -13'd374,  13'd1691,  13'd167,  13'd560,  13'd86,  -13'd398,  -13'd897,  -13'd475,  13'd2485,  13'd178,  13'd1252,  13'd1113,  -13'd1152,  13'd1004,  -13'd370,  

-13'd9,  -13'd120,  13'd689,  13'd309,  13'd208,  13'd323,  -13'd624,  13'd580,  13'd682,  13'd342,  -13'd275,  13'd863,  -13'd398,  13'd218,  -13'd62,  -13'd31,  
-13'd245,  -13'd352,  13'd630,  13'd15,  -13'd163,  -13'd240,  -13'd562,  13'd611,  13'd253,  13'd254,  -13'd546,  -13'd390,  13'd234,  13'd578,  13'd487,  -13'd111,  
13'd532,  -13'd1036,  13'd375,  -13'd201,  -13'd121,  -13'd143,  13'd340,  -13'd35,  13'd449,  -13'd26,  -13'd79,  -13'd395,  -13'd398,  13'd1074,  -13'd276,  -13'd202,  
-13'd659,  -13'd893,  -13'd584,  -13'd582,  -13'd345,  13'd503,  13'd682,  13'd202,  -13'd61,  13'd234,  13'd79,  -13'd232,  -13'd133,  13'd1134,  -13'd361,  -13'd437,  
13'd1130,  13'd1007,  -13'd125,  -13'd187,  13'd624,  13'd220,  13'd315,  -13'd81,  13'd495,  13'd265,  13'd25,  13'd171,  -13'd274,  -13'd37,  -13'd451,  13'd22,  
-13'd447,  -13'd128,  -13'd61,  13'd669,  13'd1240,  13'd475,  -13'd732,  13'd396,  -13'd1,  -13'd20,  13'd32,  13'd281,  13'd397,  13'd988,  -13'd237,  13'd843,  
-13'd885,  13'd764,  13'd219,  13'd132,  -13'd518,  -13'd513,  13'd347,  -13'd87,  -13'd377,  -13'd25,  -13'd673,  13'd130,  13'd308,  -13'd110,  13'd769,  13'd179,  
13'd229,  -13'd248,  13'd201,  13'd326,  -13'd118,  -13'd14,  13'd122,  -13'd33,  13'd51,  -13'd498,  13'd700,  -13'd5,  -13'd365,  13'd163,  -13'd25,  13'd31,  
13'd750,  -13'd393,  13'd427,  13'd376,  -13'd108,  -13'd250,  13'd804,  13'd620,  13'd134,  -13'd138,  13'd8,  -13'd103,  13'd577,  13'd209,  -13'd394,  -13'd507,  
13'd1386,  -13'd56,  -13'd824,  -13'd1,  -13'd504,  -13'd322,  13'd62,  -13'd60,  -13'd113,  -13'd755,  13'd203,  -13'd365,  13'd311,  -13'd116,  -13'd444,  13'd410,  
-13'd404,  13'd730,  -13'd869,  -13'd364,  -13'd202,  -13'd92,  -13'd403,  13'd464,  -13'd281,  13'd496,  13'd517,  -13'd1,  13'd521,  13'd154,  13'd74,  13'd15,  
-13'd134,  13'd462,  13'd161,  13'd90,  -13'd291,  13'd211,  13'd224,  -13'd333,  -13'd472,  -13'd634,  13'd389,  -13'd49,  13'd689,  13'd31,  13'd256,  13'd741,  
-13'd314,  -13'd536,  13'd303,  13'd196,  -13'd31,  13'd193,  13'd439,  13'd601,  -13'd185,  -13'd291,  13'd102,  13'd215,  13'd966,  -13'd298,  13'd345,  -13'd52,  
13'd343,  13'd8,  13'd410,  13'd600,  13'd172,  -13'd508,  13'd582,  13'd385,  13'd67,  13'd180,  13'd550,  -13'd152,  13'd391,  -13'd924,  -13'd346,  -13'd461,  
-13'd891,  -13'd285,  -13'd665,  -13'd664,  13'd311,  -13'd81,  13'd271,  13'd2,  -13'd899,  13'd143,  13'd495,  -13'd240,  13'd114,  -13'd683,  -13'd280,  13'd103,  
-13'd82,  13'd268,  -13'd553,  -13'd415,  13'd914,  13'd89,  -13'd253,  13'd184,  13'd363,  13'd164,  13'd950,  13'd172,  -13'd758,  -13'd130,  -13'd644,  -13'd129,  
-13'd209,  13'd437,  -13'd100,  -13'd699,  13'd382,  -13'd77,  13'd1206,  -13'd106,  -13'd134,  13'd328,  13'd290,  -13'd146,  13'd204,  -13'd404,  -13'd84,  13'd451,  
-13'd8,  13'd227,  13'd141,  13'd76,  -13'd620,  13'd417,  13'd271,  -13'd140,  13'd739,  13'd319,  -13'd487,  -13'd814,  -13'd21,  13'd170,  -13'd246,  13'd87,  
13'd140,  -13'd470,  13'd114,  13'd315,  -13'd854,  13'd395,  -13'd23,  -13'd124,  13'd109,  13'd292,  13'd937,  13'd54,  -13'd273,  13'd673,  -13'd78,  13'd240,  
-13'd218,  -13'd726,  13'd345,  -13'd57,  13'd319,  13'd40,  13'd73,  13'd111,  13'd233,  -13'd591,  13'd101,  13'd327,  -13'd215,  -13'd97,  -13'd379,  13'd247,  
-13'd510,  -13'd682,  -13'd574,  13'd257,  13'd174,  -13'd89,  -13'd128,  -13'd274,  13'd599,  13'd105,  -13'd62,  -13'd213,  13'd203,  -13'd828,  13'd54,  -13'd40,  
-13'd406,  -13'd128,  -13'd250,  -13'd305,  -13'd430,  -13'd274,  13'd555,  13'd535,  13'd1079,  13'd359,  13'd384,  13'd125,  13'd77,  13'd764,  -13'd325,  13'd686,  
13'd844,  13'd132,  13'd362,  13'd470,  13'd183,  -13'd383,  13'd806,  -13'd259,  13'd112,  13'd1027,  -13'd150,  13'd115,  -13'd299,  13'd1198,  13'd139,  13'd79,  
13'd670,  13'd163,  13'd294,  -13'd299,  13'd5,  13'd220,  -13'd71,  -13'd270,  -13'd420,  -13'd74,  13'd442,  -13'd150,  -13'd233,  13'd378,  13'd89,  13'd186,  
13'd761,  -13'd160,  13'd372,  13'd559,  -13'd34,  13'd22,  13'd344,  13'd156,  -13'd1007,  -13'd1154,  13'd349,  -13'd230,  -13'd70,  13'd402,  -13'd166,  13'd228,  

13'd669,  13'd136,  13'd400,  -13'd45,  13'd120,  -13'd130,  -13'd680,  13'd13,  13'd279,  13'd526,  -13'd989,  13'd181,  -13'd264,  -13'd748,  13'd604,  13'd994,  
-13'd63,  13'd279,  13'd1247,  13'd118,  13'd200,  -13'd477,  13'd408,  13'd876,  -13'd1084,  13'd228,  -13'd888,  -13'd15,  -13'd1379,  13'd807,  -13'd615,  13'd4,  
-13'd366,  -13'd961,  13'd632,  -13'd571,  -13'd875,  -13'd388,  13'd839,  13'd327,  13'd72,  13'd33,  -13'd901,  -13'd153,  -13'd556,  13'd995,  13'd163,  -13'd1160,  
-13'd1003,  13'd689,  13'd360,  -13'd417,  -13'd1006,  -13'd258,  13'd446,  -13'd59,  13'd136,  13'd131,  -13'd17,  -13'd554,  -13'd710,  -13'd361,  -13'd656,  -13'd1351,  
-13'd697,  13'd111,  -13'd415,  -13'd482,  -13'd1018,  -13'd783,  -13'd887,  -13'd682,  -13'd801,  -13'd269,  -13'd455,  -13'd622,  -13'd1261,  -13'd938,  13'd165,  -13'd620,  
-13'd420,  -13'd312,  -13'd806,  13'd517,  13'd430,  13'd786,  13'd540,  -13'd282,  -13'd330,  -13'd281,  -13'd212,  13'd331,  13'd429,  -13'd41,  -13'd754,  -13'd15,  
13'd388,  13'd569,  13'd1624,  13'd61,  13'd0,  13'd959,  13'd1130,  13'd919,  -13'd430,  13'd156,  -13'd181,  13'd532,  13'd164,  13'd805,  13'd189,  -13'd42,  
-13'd1303,  13'd736,  13'd129,  13'd112,  -13'd485,  13'd590,  13'd1002,  13'd1151,  13'd169,  13'd791,  -13'd178,  -13'd750,  13'd503,  -13'd137,  -13'd129,  -13'd1192,  
13'd702,  -13'd765,  13'd654,  -13'd41,  -13'd138,  -13'd629,  -13'd948,  -13'd246,  -13'd182,  13'd881,  -13'd516,  13'd457,  13'd298,  13'd21,  13'd264,  13'd154,  
13'd635,  13'd54,  13'd138,  -13'd271,  13'd362,  13'd406,  -13'd455,  -13'd626,  13'd48,  13'd802,  -13'd1054,  13'd689,  -13'd798,  -13'd668,  13'd120,  -13'd253,  
-13'd416,  13'd179,  -13'd52,  13'd101,  13'd504,  13'd548,  13'd509,  -13'd604,  13'd21,  13'd174,  13'd62,  13'd339,  13'd103,  13'd557,  13'd396,  13'd643,  
-13'd702,  13'd37,  -13'd166,  -13'd875,  13'd401,  -13'd55,  13'd1471,  -13'd283,  -13'd501,  -13'd235,  -13'd296,  -13'd356,  -13'd182,  13'd384,  13'd637,  -13'd577,  
-13'd340,  13'd510,  13'd231,  13'd790,  13'd195,  -13'd83,  -13'd202,  -13'd571,  13'd405,  -13'd611,  13'd823,  -13'd138,  13'd196,  13'd246,  13'd105,  13'd518,  
13'd231,  13'd367,  13'd620,  -13'd3,  13'd38,  -13'd422,  -13'd440,  -13'd364,  13'd35,  13'd330,  13'd511,  -13'd591,  13'd305,  13'd541,  13'd677,  -13'd62,  
13'd149,  -13'd430,  13'd273,  13'd603,  13'd216,  -13'd375,  13'd442,  -13'd453,  13'd99,  -13'd155,  13'd189,  13'd45,  13'd497,  -13'd847,  13'd338,  13'd172,  
-13'd302,  -13'd50,  13'd483,  -13'd456,  -13'd350,  13'd166,  13'd633,  13'd362,  13'd186,  -13'd237,  13'd550,  -13'd366,  -13'd238,  -13'd296,  13'd102,  -13'd686,  
-13'd447,  -13'd2,  13'd49,  -13'd310,  13'd714,  13'd80,  13'd169,  -13'd445,  -13'd555,  13'd164,  -13'd680,  13'd452,  -13'd312,  -13'd134,  13'd125,  13'd341,  
13'd246,  -13'd36,  13'd546,  -13'd814,  13'd443,  13'd0,  13'd202,  -13'd262,  13'd326,  -13'd30,  -13'd840,  13'd157,  -13'd833,  13'd811,  13'd913,  13'd91,  
13'd1150,  -13'd500,  13'd647,  -13'd335,  -13'd686,  -13'd476,  -13'd104,  -13'd623,  13'd499,  13'd422,  13'd107,  13'd434,  -13'd27,  13'd212,  13'd457,  13'd325,  
13'd176,  13'd814,  13'd1138,  13'd316,  -13'd3,  13'd1000,  13'd332,  -13'd247,  13'd845,  13'd163,  -13'd405,  13'd167,  13'd217,  13'd173,  -13'd129,  -13'd189,  
13'd279,  -13'd540,  13'd367,  -13'd1498,  -13'd401,  -13'd849,  -13'd86,  -13'd125,  -13'd1010,  -13'd27,  -13'd784,  -13'd383,  -13'd682,  -13'd40,  -13'd298,  -13'd746,  
-13'd82,  13'd111,  -13'd666,  -13'd628,  -13'd210,  -13'd389,  -13'd406,  -13'd489,  -13'd407,  -13'd264,  -13'd1060,  -13'd96,  -13'd736,  -13'd478,  -13'd141,  -13'd839,  
13'd846,  -13'd331,  13'd347,  -13'd753,  -13'd957,  13'd837,  13'd35,  13'd299,  -13'd345,  -13'd549,  -13'd425,  -13'd597,  13'd178,  13'd635,  13'd406,  13'd148,  
13'd363,  13'd273,  13'd326,  -13'd54,  -13'd265,  -13'd7,  13'd317,  13'd752,  -13'd581,  -13'd137,  -13'd421,  -13'd322,  -13'd439,  13'd76,  13'd971,  -13'd261,  
-13'd323,  13'd349,  13'd257,  -13'd413,  13'd492,  13'd374,  13'd475,  13'd1292,  -13'd237,  13'd38,  -13'd658,  -13'd648,  13'd6,  13'd611,  -13'd48,  13'd404,  

13'd11,  13'd155,  13'd241,  -13'd259,  -13'd676,  -13'd303,  -13'd485,  13'd101,  -13'd765,  13'd442,  -13'd87,  13'd628,  13'd431,  13'd313,  -13'd54,  -13'd154,  
-13'd294,  -13'd59,  -13'd627,  -13'd303,  13'd322,  13'd583,  -13'd203,  -13'd125,  -13'd332,  -13'd587,  13'd705,  13'd369,  -13'd502,  -13'd659,  -13'd785,  13'd327,  
-13'd20,  -13'd236,  -13'd299,  13'd609,  -13'd539,  -13'd261,  13'd176,  13'd576,  13'd23,  13'd202,  -13'd31,  -13'd59,  -13'd3,  13'd191,  13'd660,  -13'd106,  
-13'd53,  -13'd294,  13'd237,  -13'd705,  13'd78,  13'd426,  -13'd302,  13'd162,  -13'd167,  -13'd367,  13'd480,  13'd24,  13'd212,  -13'd719,  13'd295,  -13'd641,  
-13'd179,  -13'd273,  -13'd704,  -13'd651,  -13'd3,  -13'd282,  13'd303,  13'd162,  -13'd313,  -13'd913,  13'd238,  13'd102,  -13'd471,  -13'd631,  13'd370,  -13'd263,  
-13'd152,  -13'd405,  13'd143,  13'd472,  -13'd253,  -13'd95,  -13'd313,  -13'd575,  -13'd122,  -13'd357,  -13'd679,  -13'd172,  13'd271,  -13'd337,  13'd44,  13'd51,  
13'd185,  13'd673,  13'd302,  -13'd474,  -13'd486,  13'd598,  13'd45,  -13'd195,  -13'd543,  13'd496,  -13'd274,  -13'd151,  -13'd599,  13'd532,  13'd42,  13'd195,  
13'd471,  13'd452,  -13'd698,  13'd20,  13'd146,  -13'd184,  -13'd286,  -13'd278,  -13'd235,  13'd130,  -13'd596,  -13'd555,  -13'd16,  -13'd554,  -13'd476,  13'd476,  
13'd56,  13'd262,  13'd236,  -13'd641,  -13'd264,  -13'd210,  13'd447,  -13'd226,  13'd493,  -13'd901,  -13'd111,  -13'd159,  13'd21,  -13'd243,  -13'd63,  -13'd819,  
-13'd98,  -13'd2,  13'd752,  13'd132,  -13'd188,  -13'd550,  -13'd392,  -13'd278,  -13'd65,  13'd32,  -13'd233,  13'd338,  13'd48,  13'd315,  13'd413,  13'd268,  
13'd253,  13'd283,  13'd530,  13'd130,  13'd62,  -13'd236,  13'd292,  13'd388,  -13'd601,  -13'd421,  13'd217,  13'd542,  -13'd681,  -13'd751,  13'd289,  -13'd615,  
13'd320,  13'd126,  -13'd316,  -13'd533,  -13'd297,  13'd448,  -13'd313,  -13'd401,  -13'd44,  13'd223,  -13'd60,  13'd202,  13'd369,  -13'd819,  -13'd138,  -13'd207,  
-13'd359,  13'd229,  -13'd253,  -13'd197,  13'd109,  -13'd331,  13'd115,  -13'd386,  13'd62,  -13'd339,  -13'd446,  -13'd694,  -13'd741,  13'd342,  -13'd38,  13'd112,  
-13'd171,  -13'd752,  -13'd85,  -13'd265,  -13'd418,  -13'd482,  -13'd121,  -13'd82,  -13'd41,  -13'd215,  13'd57,  13'd46,  13'd180,  -13'd309,  -13'd237,  13'd339,  
-13'd52,  -13'd313,  -13'd519,  -13'd6,  -13'd111,  -13'd648,  -13'd315,  13'd131,  -13'd108,  13'd140,  -13'd6,  -13'd681,  13'd170,  -13'd289,  -13'd116,  13'd398,  
-13'd437,  13'd176,  -13'd376,  13'd660,  -13'd19,  -13'd411,  -13'd143,  -13'd163,  -13'd267,  13'd81,  13'd229,  -13'd62,  -13'd733,  -13'd404,  -13'd178,  13'd573,  
13'd37,  -13'd208,  -13'd356,  -13'd589,  -13'd238,  -13'd367,  13'd87,  -13'd237,  -13'd107,  -13'd179,  -13'd39,  -13'd490,  13'd130,  13'd226,  -13'd371,  -13'd407,  
-13'd597,  13'd163,  13'd159,  13'd444,  -13'd3,  -13'd187,  -13'd687,  13'd93,  13'd236,  13'd398,  -13'd761,  -13'd842,  -13'd544,  13'd336,  -13'd363,  -13'd271,  
-13'd533,  -13'd175,  13'd471,  -13'd224,  13'd161,  13'd20,  13'd378,  -13'd311,  -13'd392,  -13'd265,  -13'd117,  -13'd674,  -13'd429,  -13'd420,  13'd5,  13'd222,  
13'd71,  13'd93,  -13'd363,  -13'd476,  -13'd137,  13'd621,  -13'd125,  -13'd211,  13'd324,  -13'd644,  13'd53,  -13'd324,  13'd63,  -13'd206,  13'd372,  -13'd164,  
-13'd774,  13'd42,  13'd164,  -13'd477,  -13'd240,  13'd408,  -13'd12,  13'd223,  -13'd384,  -13'd411,  -13'd605,  13'd58,  -13'd397,  -13'd65,  -13'd393,  13'd3,  
-13'd821,  13'd732,  -13'd209,  -13'd433,  -13'd231,  13'd415,  13'd124,  -13'd334,  -13'd54,  -13'd124,  13'd134,  -13'd7,  -13'd482,  -13'd88,  -13'd251,  -13'd234,  
13'd316,  -13'd333,  13'd87,  -13'd149,  13'd48,  -13'd49,  -13'd96,  -13'd158,  -13'd272,  13'd56,  13'd111,  -13'd441,  -13'd812,  -13'd44,  -13'd163,  -13'd532,  
-13'd352,  -13'd144,  13'd22,  -13'd386,  -13'd79,  13'd192,  13'd148,  -13'd161,  13'd633,  -13'd71,  -13'd378,  13'd691,  13'd133,  13'd64,  -13'd447,  -13'd427,  
-13'd101,  13'd486,  13'd360,  -13'd220,  -13'd59,  13'd56,  -13'd299,  13'd300,  -13'd206,  -13'd414,  -13'd612,  13'd398,  -13'd760,  -13'd877,  -13'd209,  -13'd46,  

-13'd46,  13'd213,  -13'd629,  13'd317,  -13'd830,  -13'd362,  -13'd567,  -13'd441,  13'd75,  -13'd436,  13'd642,  13'd79,  -13'd391,  -13'd830,  -13'd406,  -13'd605,  
-13'd125,  -13'd708,  -13'd439,  13'd100,  -13'd10,  -13'd597,  -13'd649,  13'd588,  13'd479,  13'd334,  -13'd48,  13'd247,  -13'd605,  -13'd749,  13'd272,  -13'd170,  
13'd186,  -13'd684,  -13'd204,  13'd95,  -13'd180,  13'd14,  -13'd975,  -13'd274,  -13'd593,  13'd1053,  13'd374,  -13'd439,  13'd367,  -13'd1860,  -13'd137,  13'd21,  
-13'd602,  -13'd1617,  -13'd615,  13'd784,  13'd497,  13'd458,  -13'd619,  13'd185,  13'd734,  13'd637,  -13'd399,  -13'd328,  -13'd103,  -13'd983,  -13'd526,  13'd135,  
-13'd1533,  -13'd838,  13'd335,  13'd168,  -13'd39,  13'd166,  13'd72,  13'd253,  -13'd386,  13'd15,  -13'd769,  -13'd653,  13'd313,  -13'd217,  13'd101,  -13'd1211,  
13'd191,  13'd141,  13'd15,  13'd142,  -13'd111,  13'd793,  13'd120,  13'd72,  -13'd155,  -13'd269,  13'd536,  13'd4,  -13'd937,  -13'd296,  -13'd351,  13'd344,  
13'd599,  13'd851,  -13'd74,  13'd156,  -13'd22,  -13'd465,  13'd46,  -13'd93,  13'd531,  13'd56,  -13'd430,  -13'd15,  13'd167,  -13'd683,  -13'd212,  13'd484,  
13'd78,  -13'd194,  -13'd879,  -13'd483,  -13'd170,  13'd838,  -13'd50,  -13'd608,  -13'd83,  -13'd200,  13'd79,  13'd579,  13'd182,  -13'd349,  13'd174,  -13'd0,  
-13'd302,  13'd635,  13'd343,  13'd767,  -13'd363,  -13'd415,  13'd368,  13'd527,  13'd1091,  13'd929,  13'd356,  13'd288,  13'd31,  13'd75,  13'd54,  -13'd18,  
-13'd1358,  -13'd943,  -13'd596,  13'd125,  -13'd395,  -13'd557,  13'd270,  13'd32,  13'd383,  -13'd746,  13'd275,  -13'd566,  -13'd482,  13'd70,  -13'd314,  -13'd307,  
13'd0,  13'd155,  -13'd9,  -13'd96,  13'd25,  13'd719,  13'd464,  13'd397,  -13'd75,  13'd247,  -13'd931,  13'd77,  13'd536,  13'd435,  -13'd8,  -13'd66,  
-13'd230,  13'd89,  13'd342,  13'd78,  -13'd348,  -13'd349,  13'd131,  13'd238,  13'd128,  -13'd282,  -13'd174,  13'd434,  13'd176,  -13'd632,  13'd322,  -13'd213,  
-13'd173,  13'd491,  -13'd212,  -13'd329,  13'd100,  -13'd574,  -13'd530,  -13'd338,  -13'd693,  13'd120,  13'd431,  -13'd267,  13'd344,  -13'd602,  -13'd70,  13'd300,  
13'd911,  -13'd178,  -13'd40,  -13'd198,  13'd449,  13'd547,  13'd243,  -13'd268,  -13'd131,  -13'd660,  13'd601,  13'd287,  -13'd452,  13'd326,  -13'd101,  13'd144,  
13'd411,  -13'd355,  13'd571,  -13'd51,  13'd247,  -13'd20,  13'd478,  13'd691,  13'd259,  -13'd919,  13'd420,  13'd667,  13'd63,  13'd574,  13'd179,  13'd71,  
13'd151,  -13'd53,  13'd144,  -13'd188,  13'd747,  13'd462,  -13'd231,  13'd9,  -13'd438,  -13'd93,  -13'd305,  13'd224,  13'd86,  13'd790,  -13'd12,  -13'd570,  
13'd39,  -13'd86,  -13'd691,  -13'd35,  -13'd184,  -13'd198,  -13'd531,  13'd552,  13'd4,  -13'd862,  13'd414,  -13'd548,  13'd7,  13'd261,  13'd257,  13'd575,  
-13'd527,  13'd666,  -13'd151,  -13'd514,  13'd96,  -13'd67,  13'd81,  13'd581,  -13'd386,  13'd28,  13'd537,  -13'd257,  -13'd463,  13'd196,  -13'd703,  13'd209,  
13'd794,  13'd789,  13'd411,  -13'd510,  -13'd562,  13'd173,  -13'd31,  -13'd481,  -13'd305,  13'd418,  13'd267,  13'd158,  13'd313,  13'd209,  13'd418,  -13'd347,  
13'd348,  13'd671,  -13'd681,  13'd37,  13'd225,  13'd190,  -13'd232,  13'd493,  -13'd662,  -13'd438,  -13'd268,  -13'd598,  -13'd16,  -13'd79,  13'd518,  13'd136,  
-13'd49,  13'd575,  -13'd94,  -13'd410,  13'd287,  -13'd256,  -13'd646,  -13'd731,  13'd311,  13'd312,  -13'd25,  13'd6,  -13'd914,  -13'd190,  -13'd62,  -13'd331,  
-13'd511,  -13'd795,  13'd655,  13'd163,  -13'd149,  -13'd406,  13'd229,  -13'd251,  13'd337,  13'd122,  13'd140,  -13'd72,  -13'd738,  -13'd420,  -13'd41,  -13'd7,  
-13'd690,  -13'd193,  13'd292,  -13'd280,  13'd86,  13'd392,  13'd747,  -13'd536,  13'd1031,  13'd818,  -13'd252,  -13'd390,  -13'd592,  13'd1076,  13'd347,  13'd122,  
-13'd381,  -13'd159,  -13'd291,  -13'd698,  13'd79,  13'd546,  -13'd601,  13'd83,  13'd281,  13'd239,  13'd74,  13'd3,  13'd266,  13'd397,  13'd117,  -13'd564,  
-13'd527,  -13'd498,  13'd184,  13'd639,  -13'd811,  -13'd95,  -13'd408,  13'd21,  13'd66,  13'd169,  -13'd507,  -13'd253,  13'd52,  -13'd897,  13'd400,  -13'd556,  

-13'd121,  -13'd34,  -13'd539,  13'd210,  13'd163,  -13'd283,  -13'd110,  13'd208,  -13'd610,  -13'd477,  -13'd617,  13'd235,  -13'd233,  13'd66,  13'd236,  -13'd1028,  
13'd84,  13'd721,  -13'd558,  -13'd256,  13'd708,  -13'd12,  -13'd645,  -13'd276,  13'd209,  13'd266,  -13'd319,  13'd266,  -13'd200,  -13'd491,  13'd123,  -13'd180,  
-13'd188,  13'd627,  -13'd752,  -13'd198,  13'd318,  13'd219,  13'd761,  -13'd283,  -13'd582,  13'd297,  13'd262,  13'd437,  -13'd91,  -13'd560,  -13'd253,  13'd297,  
-13'd698,  -13'd189,  13'd287,  -13'd601,  13'd644,  -13'd619,  13'd69,  -13'd689,  13'd366,  -13'd415,  -13'd694,  13'd659,  13'd143,  13'd360,  -13'd382,  13'd549,  
-13'd598,  -13'd963,  -13'd345,  -13'd599,  -13'd410,  -13'd90,  -13'd365,  -13'd129,  -13'd48,  -13'd446,  -13'd175,  -13'd709,  -13'd284,  13'd133,  -13'd504,  -13'd233,  
13'd126,  13'd161,  -13'd85,  13'd417,  -13'd106,  13'd108,  13'd35,  -13'd103,  13'd824,  -13'd242,  -13'd59,  13'd109,  13'd226,  13'd426,  -13'd523,  -13'd390,  
13'd440,  13'd3,  -13'd153,  -13'd507,  -13'd625,  13'd135,  -13'd221,  13'd395,  -13'd507,  -13'd228,  -13'd364,  -13'd271,  13'd479,  -13'd239,  -13'd426,  13'd527,  
13'd779,  -13'd0,  -13'd95,  -13'd132,  -13'd473,  -13'd267,  13'd254,  13'd774,  -13'd377,  -13'd265,  -13'd419,  13'd562,  13'd452,  13'd258,  13'd819,  13'd123,  
-13'd16,  -13'd93,  13'd56,  -13'd130,  13'd21,  13'd175,  13'd1067,  -13'd409,  13'd205,  -13'd261,  -13'd25,  13'd962,  13'd194,  13'd1409,  13'd119,  -13'd214,  
-13'd576,  13'd21,  -13'd271,  -13'd223,  13'd116,  13'd130,  13'd439,  13'd472,  -13'd199,  13'd296,  -13'd64,  -13'd809,  -13'd114,  13'd331,  -13'd303,  -13'd887,  
-13'd89,  -13'd4,  -13'd169,  -13'd98,  13'd717,  13'd153,  -13'd126,  -13'd245,  -13'd119,  13'd148,  -13'd901,  -13'd229,  -13'd616,  13'd571,  -13'd566,  -13'd267,  
13'd308,  13'd114,  13'd905,  13'd442,  13'd621,  -13'd44,  -13'd548,  -13'd329,  -13'd201,  -13'd700,  13'd116,  13'd570,  13'd79,  -13'd430,  13'd214,  -13'd228,  
13'd234,  13'd277,  13'd198,  -13'd514,  -13'd706,  13'd819,  -13'd416,  13'd706,  13'd238,  -13'd469,  13'd937,  13'd217,  13'd271,  13'd197,  -13'd577,  13'd709,  
-13'd553,  -13'd2,  13'd444,  13'd593,  -13'd698,  -13'd338,  13'd364,  13'd189,  13'd393,  -13'd234,  13'd365,  -13'd292,  13'd238,  13'd390,  13'd363,  -13'd286,  
13'd253,  -13'd446,  -13'd43,  13'd16,  13'd72,  -13'd528,  -13'd396,  -13'd214,  13'd260,  -13'd598,  -13'd38,  -13'd977,  13'd449,  13'd490,  -13'd262,  -13'd712,  
-13'd411,  -13'd204,  -13'd704,  13'd138,  -13'd641,  13'd388,  -13'd169,  -13'd363,  -13'd126,  13'd322,  -13'd166,  -13'd673,  -13'd122,  13'd39,  -13'd524,  13'd274,  
-13'd88,  13'd54,  -13'd391,  13'd450,  -13'd137,  -13'd67,  -13'd371,  13'd726,  13'd309,  -13'd675,  13'd886,  -13'd436,  13'd71,  13'd11,  13'd99,  13'd30,  
13'd275,  -13'd194,  13'd793,  -13'd208,  13'd596,  -13'd575,  -13'd234,  -13'd117,  13'd667,  13'd716,  13'd318,  13'd216,  13'd396,  -13'd32,  -13'd813,  -13'd267,  
13'd466,  -13'd249,  13'd115,  -13'd164,  -13'd513,  13'd243,  -13'd15,  13'd227,  13'd468,  13'd15,  13'd129,  -13'd212,  -13'd187,  13'd637,  13'd64,  -13'd687,  
13'd305,  -13'd700,  -13'd1096,  -13'd620,  -13'd597,  -13'd574,  -13'd147,  -13'd591,  -13'd932,  13'd675,  -13'd391,  -13'd176,  13'd86,  13'd226,  -13'd62,  -13'd791,  
13'd107,  13'd30,  13'd59,  -13'd218,  13'd569,  -13'd187,  13'd599,  -13'd702,  -13'd776,  13'd399,  13'd685,  13'd238,  -13'd429,  13'd334,  -13'd19,  13'd608,  
-13'd84,  13'd103,  -13'd405,  13'd216,  13'd89,  -13'd346,  13'd730,  -13'd14,  13'd1083,  -13'd0,  13'd338,  -13'd446,  -13'd754,  -13'd131,  13'd82,  13'd475,  
-13'd128,  13'd101,  13'd383,  -13'd227,  13'd435,  -13'd301,  -13'd692,  -13'd123,  13'd104,  -13'd541,  -13'd928,  -13'd134,  13'd128,  13'd1065,  13'd118,  13'd129,  
-13'd194,  13'd75,  -13'd74,  13'd207,  -13'd278,  13'd339,  -13'd535,  -13'd456,  -13'd161,  13'd567,  -13'd59,  -13'd65,  -13'd752,  -13'd21,  13'd789,  13'd658,  
-13'd959,  13'd208,  13'd681,  13'd80,  13'd69,  13'd726,  13'd563,  -13'd712,  13'd46,  13'd1465,  13'd498,  -13'd643,  -13'd147,  -13'd584,  13'd378,  -13'd296,  

-13'd742,  13'd411,  -13'd201,  13'd631,  -13'd103,  13'd215,  -13'd91,  -13'd483,  13'd472,  -13'd10,  13'd106,  13'd473,  13'd200,  13'd153,  13'd40,  13'd57,  
-13'd381,  13'd615,  13'd97,  13'd687,  -13'd72,  -13'd96,  -13'd406,  13'd828,  -13'd663,  13'd104,  -13'd410,  13'd682,  -13'd149,  13'd501,  -13'd190,  13'd459,  
-13'd379,  -13'd897,  13'd742,  -13'd520,  13'd164,  13'd107,  13'd306,  -13'd232,  13'd875,  13'd45,  -13'd180,  -13'd564,  13'd381,  13'd1186,  13'd266,  -13'd175,  
-13'd384,  -13'd909,  -13'd549,  13'd16,  -13'd456,  13'd177,  13'd159,  -13'd32,  -13'd455,  -13'd68,  13'd496,  13'd653,  -13'd408,  -13'd543,  -13'd234,  -13'd277,  
-13'd264,  -13'd574,  -13'd480,  -13'd141,  -13'd368,  -13'd84,  13'd766,  -13'd69,  -13'd685,  -13'd776,  13'd54,  -13'd269,  -13'd190,  13'd329,  13'd21,  13'd218,  
-13'd396,  13'd257,  -13'd275,  -13'd316,  -13'd330,  13'd41,  -13'd370,  13'd33,  -13'd787,  -13'd307,  13'd356,  13'd47,  13'd292,  13'd685,  -13'd129,  13'd61,  
13'd468,  -13'd542,  13'd263,  13'd32,  -13'd86,  -13'd232,  13'd216,  -13'd351,  -13'd625,  -13'd23,  -13'd19,  13'd91,  -13'd538,  -13'd50,  13'd191,  13'd400,  
13'd23,  -13'd688,  -13'd139,  13'd29,  -13'd265,  -13'd263,  -13'd135,  13'd510,  13'd637,  -13'd492,  13'd140,  -13'd113,  -13'd8,  -13'd111,  13'd523,  13'd422,  
-13'd188,  -13'd914,  13'd2,  13'd125,  -13'd485,  -13'd160,  -13'd68,  13'd268,  -13'd109,  -13'd103,  13'd22,  -13'd173,  -13'd73,  -13'd108,  13'd188,  -13'd634,  
-13'd584,  13'd166,  -13'd740,  -13'd120,  -13'd913,  13'd806,  -13'd431,  13'd196,  13'd261,  -13'd325,  13'd319,  -13'd307,  13'd240,  -13'd62,  -13'd150,  13'd712,  
-13'd283,  -13'd246,  13'd118,  13'd101,  -13'd701,  -13'd789,  -13'd919,  13'd30,  13'd320,  13'd710,  13'd58,  -13'd274,  -13'd44,  -13'd117,  -13'd51,  -13'd101,  
13'd421,  -13'd606,  13'd497,  13'd31,  -13'd1005,  13'd75,  -13'd1454,  13'd207,  -13'd1006,  13'd1087,  -13'd112,  13'd375,  -13'd233,  -13'd197,  13'd340,  13'd707,  
-13'd407,  -13'd425,  -13'd343,  -13'd209,  13'd415,  -13'd332,  -13'd763,  -13'd205,  -13'd1041,  -13'd183,  -13'd195,  -13'd136,  13'd221,  13'd263,  13'd539,  13'd410,  
-13'd130,  13'd311,  -13'd623,  -13'd73,  13'd226,  -13'd684,  -13'd314,  13'd215,  -13'd378,  -13'd617,  13'd37,  13'd435,  -13'd500,  -13'd532,  -13'd332,  -13'd38,  
-13'd1844,  -13'd932,  13'd82,  -13'd314,  13'd536,  -13'd382,  -13'd640,  -13'd156,  13'd11,  13'd817,  -13'd366,  13'd325,  -13'd780,  -13'd312,  -13'd89,  -13'd882,  
-13'd1149,  -13'd1006,  -13'd174,  13'd861,  -13'd148,  -13'd207,  -13'd1770,  13'd433,  13'd407,  13'd166,  13'd90,  -13'd383,  13'd78,  -13'd371,  -13'd116,  -13'd548,  
-13'd851,  -13'd661,  13'd971,  -13'd474,  13'd369,  -13'd255,  -13'd752,  -13'd411,  -13'd353,  13'd723,  13'd476,  13'd177,  -13'd102,  -13'd279,  -13'd540,  -13'd158,  
13'd326,  -13'd599,  13'd281,  13'd89,  -13'd362,  13'd323,  13'd381,  13'd261,  13'd330,  13'd164,  13'd294,  13'd235,  -13'd123,  -13'd248,  13'd40,  -13'd125,  
-13'd230,  -13'd1,  -13'd366,  13'd730,  13'd314,  13'd704,  13'd168,  13'd628,  -13'd43,  -13'd465,  13'd542,  13'd553,  13'd371,  13'd459,  13'd868,  13'd781,  
-13'd250,  -13'd193,  -13'd29,  13'd454,  -13'd70,  13'd163,  13'd600,  13'd530,  13'd921,  13'd526,  -13'd115,  13'd53,  -13'd530,  13'd318,  13'd410,  13'd141,  
-13'd518,  13'd102,  -13'd754,  13'd515,  13'd87,  13'd551,  -13'd37,  13'd285,  13'd1794,  13'd565,  13'd617,  13'd814,  -13'd202,  -13'd525,  13'd380,  13'd168,  
-13'd149,  -13'd53,  -13'd235,  13'd812,  13'd393,  13'd93,  13'd2,  13'd255,  13'd446,  13'd182,  13'd234,  13'd339,  13'd755,  -13'd2154,  13'd196,  13'd555,  
13'd561,  13'd441,  -13'd565,  -13'd269,  13'd410,  13'd249,  -13'd311,  13'd446,  13'd483,  13'd376,  13'd142,  13'd61,  13'd1025,  -13'd668,  -13'd63,  -13'd38,  
13'd881,  13'd490,  -13'd252,  -13'd244,  13'd43,  13'd314,  13'd354,  13'd546,  13'd431,  -13'd74,  -13'd255,  -13'd411,  13'd581,  13'd127,  -13'd156,  13'd240,  
13'd730,  13'd1032,  13'd22,  13'd364,  -13'd482,  13'd468,  -13'd341,  13'd57,  13'd422,  -13'd311,  -13'd336,  13'd108,  13'd494,  13'd464,  13'd255,  13'd167,  

-13'd260,  13'd118,  13'd250,  13'd395,  -13'd393,  -13'd65,  -13'd91,  13'd9,  -13'd233,  13'd477,  13'd437,  -13'd380,  13'd436,  -13'd130,  -13'd66,  13'd463,  
13'd126,  13'd106,  13'd414,  -13'd334,  -13'd83,  -13'd152,  -13'd838,  -13'd495,  13'd748,  -13'd55,  -13'd310,  -13'd332,  13'd213,  -13'd430,  13'd59,  -13'd198,  
-13'd121,  13'd184,  13'd405,  -13'd443,  -13'd67,  13'd250,  -13'd375,  13'd64,  13'd88,  13'd513,  13'd221,  -13'd238,  -13'd627,  13'd158,  -13'd1,  -13'd769,  
-13'd432,  -13'd479,  -13'd304,  13'd40,  13'd401,  -13'd121,  13'd96,  -13'd273,  13'd78,  -13'd16,  -13'd66,  13'd506,  13'd5,  -13'd341,  13'd128,  -13'd777,  
13'd315,  13'd160,  -13'd426,  -13'd92,  -13'd162,  13'd95,  -13'd817,  -13'd426,  13'd310,  -13'd374,  13'd512,  -13'd51,  13'd320,  -13'd81,  13'd299,  -13'd94,  
-13'd361,  13'd436,  13'd121,  13'd20,  13'd66,  -13'd644,  -13'd524,  13'd76,  -13'd249,  13'd249,  13'd583,  -13'd313,  13'd641,  13'd64,  -13'd332,  13'd381,  
13'd699,  -13'd610,  -13'd352,  -13'd318,  -13'd341,  -13'd169,  13'd230,  13'd495,  -13'd297,  -13'd50,  -13'd702,  -13'd558,  -13'd255,  13'd326,  -13'd151,  -13'd161,  
13'd291,  -13'd265,  -13'd107,  -13'd471,  -13'd596,  -13'd207,  13'd149,  13'd218,  -13'd807,  13'd57,  -13'd624,  -13'd631,  13'd128,  -13'd383,  -13'd512,  -13'd563,  
-13'd138,  13'd157,  -13'd393,  13'd28,  -13'd917,  13'd159,  13'd184,  -13'd88,  -13'd218,  -13'd430,  13'd421,  -13'd524,  13'd46,  -13'd44,  13'd197,  13'd103,  
-13'd211,  13'd541,  -13'd499,  13'd261,  -13'd474,  -13'd221,  -13'd423,  -13'd307,  -13'd801,  -13'd17,  13'd659,  13'd313,  13'd86,  13'd39,  -13'd817,  13'd196,  
13'd194,  -13'd292,  -13'd787,  -13'd690,  13'd41,  -13'd90,  -13'd392,  -13'd494,  13'd28,  13'd243,  -13'd172,  13'd11,  -13'd680,  -13'd681,  13'd49,  13'd392,  
-13'd717,  -13'd602,  13'd510,  13'd46,  -13'd216,  -13'd589,  13'd592,  -13'd302,  13'd298,  -13'd105,  13'd520,  13'd116,  13'd329,  13'd51,  -13'd554,  -13'd642,  
-13'd205,  13'd167,  13'd72,  -13'd43,  13'd300,  13'd517,  -13'd458,  -13'd281,  -13'd465,  13'd576,  13'd86,  13'd141,  13'd77,  -13'd124,  -13'd322,  -13'd207,  
-13'd306,  -13'd121,  13'd141,  -13'd481,  -13'd317,  13'd489,  -13'd758,  13'd425,  -13'd675,  -13'd133,  13'd111,  13'd173,  13'd232,  -13'd137,  -13'd248,  -13'd28,  
-13'd132,  -13'd660,  -13'd169,  13'd90,  13'd367,  13'd402,  -13'd695,  -13'd382,  13'd300,  13'd479,  -13'd260,  -13'd39,  -13'd593,  13'd141,  13'd323,  -13'd367,  
-13'd310,  -13'd11,  13'd351,  13'd329,  13'd292,  13'd456,  13'd138,  -13'd621,  -13'd362,  -13'd303,  -13'd623,  -13'd282,  13'd208,  -13'd511,  -13'd484,  13'd637,  
13'd391,  13'd639,  13'd214,  -13'd72,  -13'd380,  -13'd181,  -13'd212,  -13'd248,  -13'd581,  -13'd324,  -13'd86,  -13'd561,  -13'd256,  13'd138,  13'd614,  13'd192,  
-13'd334,  13'd231,  -13'd46,  -13'd526,  -13'd594,  13'd351,  13'd89,  -13'd71,  13'd217,  -13'd158,  13'd29,  13'd205,  -13'd261,  13'd230,  -13'd133,  -13'd2,  
13'd263,  -13'd290,  -13'd469,  13'd206,  13'd25,  -13'd26,  -13'd176,  13'd212,  13'd699,  -13'd85,  13'd258,  -13'd328,  -13'd51,  13'd266,  -13'd15,  -13'd291,  
-13'd100,  -13'd626,  -13'd146,  -13'd190,  13'd229,  13'd224,  -13'd313,  13'd236,  -13'd100,  13'd297,  -13'd353,  13'd341,  13'd152,  -13'd358,  13'd208,  -13'd405,  
13'd14,  13'd264,  13'd779,  -13'd754,  13'd151,  -13'd265,  13'd559,  13'd45,  13'd499,  13'd243,  -13'd241,  13'd177,  13'd745,  -13'd398,  -13'd99,  -13'd150,  
-13'd411,  -13'd32,  -13'd72,  13'd256,  13'd368,  -13'd719,  13'd344,  -13'd540,  -13'd593,  13'd476,  -13'd408,  -13'd24,  13'd263,  -13'd43,  13'd49,  -13'd65,  
-13'd577,  13'd151,  -13'd119,  -13'd617,  13'd372,  -13'd615,  13'd33,  13'd510,  -13'd298,  -13'd33,  -13'd131,  13'd401,  13'd220,  -13'd14,  -13'd358,  13'd26,  
13'd167,  13'd114,  -13'd500,  13'd538,  13'd305,  -13'd306,  -13'd714,  -13'd92,  13'd612,  13'd584,  -13'd317,  13'd243,  -13'd443,  -13'd296,  13'd422,  13'd470,  
-13'd670,  13'd168,  -13'd154,  13'd332,  -13'd25,  13'd154,  13'd441,  13'd681,  -13'd23,  -13'd399,  13'd421,  13'd309,  13'd239,  13'd125,  -13'd214,  13'd354,  

13'd13,  13'd36,  -13'd811,  13'd164,  13'd338,  -13'd58,  13'd515,  13'd559,  13'd197,  -13'd652,  13'd811,  13'd286,  13'd1007,  13'd197,  13'd519,  13'd886,  
13'd37,  13'd599,  -13'd879,  13'd452,  13'd130,  13'd467,  13'd154,  13'd441,  13'd546,  13'd190,  13'd700,  -13'd206,  13'd421,  -13'd904,  13'd627,  13'd288,  
-13'd1062,  -13'd218,  13'd217,  -13'd304,  13'd475,  13'd268,  -13'd1294,  -13'd37,  -13'd679,  -13'd894,  -13'd738,  -13'd204,  13'd742,  13'd468,  13'd135,  13'd648,  
-13'd19,  -13'd685,  -13'd417,  -13'd502,  -13'd524,  -13'd328,  13'd159,  13'd176,  -13'd277,  13'd370,  13'd262,  13'd284,  -13'd740,  -13'd358,  -13'd385,  -13'd1282,  
-13'd4,  -13'd542,  -13'd104,  -13'd757,  -13'd848,  13'd80,  -13'd209,  -13'd42,  -13'd10,  -13'd111,  -13'd446,  -13'd17,  -13'd750,  13'd658,  -13'd1015,  -13'd429,  
-13'd559,  13'd546,  13'd97,  -13'd124,  13'd285,  13'd325,  13'd960,  -13'd235,  13'd91,  -13'd73,  13'd734,  13'd126,  -13'd616,  -13'd264,  -13'd726,  -13'd493,  
13'd116,  -13'd70,  -13'd71,  13'd1,  13'd412,  13'd265,  13'd3,  13'd4,  13'd428,  13'd561,  13'd410,  -13'd282,  -13'd57,  -13'd262,  13'd535,  -13'd430,  
13'd40,  13'd45,  13'd72,  -13'd149,  13'd529,  -13'd417,  -13'd629,  13'd148,  -13'd563,  -13'd55,  -13'd52,  13'd220,  -13'd358,  13'd415,  13'd7,  13'd160,  
-13'd44,  -13'd635,  -13'd864,  -13'd359,  -13'd265,  -13'd898,  -13'd312,  -13'd805,  13'd506,  -13'd565,  -13'd617,  -13'd495,  -13'd1092,  13'd502,  -13'd335,  -13'd347,  
-13'd949,  13'd239,  13'd371,  -13'd353,  -13'd389,  -13'd230,  -13'd387,  -13'd1024,  -13'd985,  13'd338,  -13'd477,  13'd111,  -13'd1128,  13'd1064,  -13'd403,  -13'd216,  
-13'd170,  -13'd94,  -13'd731,  -13'd147,  13'd147,  13'd44,  13'd731,  -13'd770,  13'd114,  -13'd472,  -13'd324,  -13'd747,  -13'd2,  13'd71,  -13'd409,  13'd118,  
-13'd285,  13'd487,  -13'd183,  -13'd40,  13'd193,  -13'd0,  -13'd215,  13'd14,  13'd1071,  13'd371,  -13'd455,  -13'd79,  13'd296,  -13'd158,  13'd537,  13'd537,  
-13'd45,  13'd329,  13'd24,  -13'd18,  -13'd263,  13'd290,  -13'd128,  -13'd60,  13'd887,  13'd451,  13'd498,  -13'd277,  13'd346,  13'd384,  -13'd395,  -13'd129,  
-13'd1154,  13'd423,  -13'd1213,  13'd1060,  13'd19,  13'd444,  13'd428,  -13'd153,  13'd993,  -13'd592,  13'd1461,  13'd239,  -13'd151,  13'd137,  -13'd345,  13'd480,  
-13'd1049,  -13'd74,  13'd823,  13'd824,  -13'd126,  -13'd151,  -13'd62,  13'd298,  -13'd202,  -13'd134,  13'd1631,  13'd79,  13'd959,  -13'd243,  13'd27,  13'd440,  
13'd1110,  13'd217,  13'd572,  -13'd486,  -13'd703,  13'd616,  -13'd394,  -13'd115,  13'd63,  13'd73,  -13'd1073,  -13'd519,  -13'd698,  13'd841,  13'd240,  -13'd941,  
13'd400,  -13'd100,  -13'd27,  -13'd192,  -13'd43,  -13'd738,  -13'd445,  -13'd288,  -13'd228,  -13'd73,  -13'd362,  -13'd196,  13'd187,  13'd467,  13'd1038,  13'd670,  
13'd303,  -13'd606,  13'd219,  -13'd750,  13'd498,  13'd43,  13'd489,  -13'd688,  13'd129,  13'd700,  13'd673,  13'd72,  -13'd177,  -13'd190,  -13'd303,  13'd198,  
-13'd12,  13'd1477,  -13'd463,  13'd344,  13'd225,  -13'd153,  13'd38,  13'd92,  13'd338,  -13'd597,  13'd799,  -13'd87,  13'd375,  13'd113,  13'd405,  13'd588,  
-13'd110,  -13'd410,  -13'd421,  13'd22,  13'd35,  -13'd747,  -13'd38,  -13'd458,  -13'd676,  13'd485,  13'd814,  -13'd665,  -13'd40,  13'd48,  13'd134,  13'd1103,  
13'd174,  13'd323,  13'd766,  13'd704,  -13'd511,  13'd329,  -13'd804,  13'd475,  -13'd930,  -13'd88,  -13'd817,  -13'd669,  -13'd526,  13'd624,  13'd140,  -13'd977,  
13'd446,  -13'd270,  -13'd423,  -13'd234,  -13'd423,  13'd14,  -13'd56,  -13'd107,  -13'd631,  -13'd273,  13'd9,  -13'd667,  13'd211,  13'd635,  13'd425,  13'd95,  
13'd260,  -13'd177,  -13'd161,  13'd324,  13'd1043,  -13'd404,  13'd738,  13'd631,  -13'd705,  -13'd878,  -13'd133,  -13'd662,  -13'd477,  -13'd367,  -13'd652,  13'd48,  
-13'd1159,  13'd639,  13'd120,  -13'd133,  13'd57,  13'd271,  -13'd453,  13'd686,  -13'd121,  13'd467,  -13'd597,  -13'd996,  -13'd585,  13'd614,  -13'd896,  13'd26,  
-13'd1153,  -13'd186,  13'd58,  13'd840,  13'd299,  -13'd133,  -13'd343,  -13'd115,  -13'd847,  13'd1404,  13'd105,  -13'd244,  -13'd205,  -13'd116,  -13'd59,  13'd227,  

-13'd609,  -13'd228,  -13'd270,  -13'd129,  13'd549,  -13'd192,  13'd253,  13'd472,  -13'd179,  13'd13,  13'd666,  -13'd838,  -13'd28,  -13'd705,  13'd625,  13'd96,  
-13'd621,  -13'd184,  -13'd5,  13'd201,  13'd265,  -13'd152,  -13'd1380,  -13'd22,  -13'd751,  13'd669,  -13'd982,  -13'd369,  13'd497,  -13'd1254,  -13'd21,  13'd14,  
-13'd194,  -13'd757,  13'd557,  13'd897,  -13'd444,  13'd215,  13'd580,  13'd685,  -13'd319,  13'd630,  13'd621,  -13'd306,  -13'd554,  -13'd936,  13'd206,  13'd711,  
13'd788,  -13'd1235,  -13'd467,  13'd385,  -13'd43,  13'd795,  13'd708,  13'd441,  13'd510,  -13'd303,  13'd146,  13'd382,  13'd622,  13'd1082,  -13'd277,  -13'd385,  
-13'd856,  -13'd28,  13'd283,  -13'd518,  13'd267,  13'd425,  13'd136,  -13'd374,  13'd804,  -13'd546,  13'd321,  13'd323,  -13'd1074,  13'd429,  -13'd91,  -13'd260,  
-13'd848,  13'd50,  -13'd682,  -13'd318,  -13'd417,  -13'd840,  -13'd1005,  -13'd44,  -13'd253,  -13'd643,  13'd716,  -13'd32,  -13'd260,  -13'd426,  -13'd12,  13'd328,  
-13'd346,  -13'd520,  -13'd852,  -13'd785,  13'd541,  13'd118,  -13'd193,  13'd196,  -13'd196,  -13'd93,  13'd628,  13'd50,  -13'd338,  -13'd558,  13'd293,  13'd262,  
13'd449,  -13'd284,  -13'd557,  13'd281,  -13'd2,  -13'd224,  -13'd51,  -13'd40,  -13'd662,  13'd536,  -13'd59,  -13'd6,  -13'd205,  -13'd857,  13'd589,  13'd547,  
13'd1040,  13'd97,  -13'd317,  -13'd81,  -13'd142,  -13'd464,  13'd718,  13'd455,  -13'd223,  13'd264,  -13'd200,  13'd77,  -13'd360,  13'd124,  13'd135,  13'd162,  
-13'd300,  13'd467,  -13'd164,  13'd545,  -13'd437,  13'd532,  13'd270,  -13'd199,  -13'd747,  -13'd21,  13'd94,  -13'd481,  13'd214,  13'd173,  -13'd337,  -13'd463,  
-13'd653,  -13'd217,  13'd124,  -13'd267,  -13'd735,  -13'd478,  13'd596,  13'd423,  13'd677,  -13'd383,  13'd521,  -13'd278,  -13'd614,  -13'd191,  13'd158,  -13'd653,  
13'd517,  -13'd481,  13'd235,  -13'd472,  -13'd937,  -13'd750,  13'd229,  -13'd206,  -13'd140,  13'd361,  -13'd677,  -13'd551,  13'd125,  13'd582,  13'd788,  -13'd541,  
13'd444,  -13'd226,  13'd597,  -13'd387,  -13'd646,  13'd151,  13'd111,  13'd152,  13'd140,  13'd134,  13'd44,  13'd374,  -13'd206,  13'd123,  -13'd312,  -13'd275,  
-13'd340,  -13'd72,  -13'd108,  13'd338,  13'd174,  13'd291,  13'd207,  13'd470,  13'd258,  13'd443,  13'd86,  13'd568,  -13'd159,  -13'd307,  13'd37,  13'd448,  
-13'd297,  -13'd29,  13'd184,  13'd157,  -13'd191,  -13'd253,  13'd242,  -13'd100,  13'd137,  13'd595,  13'd186,  -13'd391,  -13'd35,  -13'd128,  -13'd104,  -13'd434,  
-13'd692,  -13'd674,  13'd408,  13'd851,  -13'd44,  13'd607,  -13'd433,  13'd491,  13'd385,  13'd181,  13'd398,  -13'd180,  -13'd379,  13'd74,  13'd133,  13'd223,  
-13'd990,  -13'd279,  -13'd193,  13'd168,  13'd2,  -13'd425,  13'd459,  -13'd647,  -13'd411,  13'd863,  13'd626,  -13'd319,  -13'd427,  -13'd70,  13'd641,  -13'd215,  
-13'd105,  13'd422,  13'd214,  13'd271,  -13'd59,  13'd289,  13'd152,  13'd265,  -13'd244,  -13'd503,  -13'd527,  -13'd51,  -13'd13,  13'd178,  -13'd122,  -13'd540,  
13'd2,  -13'd92,  13'd627,  13'd732,  -13'd843,  -13'd283,  -13'd16,  -13'd324,  -13'd777,  -13'd490,  -13'd161,  13'd176,  13'd268,  -13'd29,  13'd75,  13'd646,  
13'd19,  13'd168,  13'd148,  13'd213,  -13'd372,  -13'd193,  13'd433,  13'd52,  -13'd469,  -13'd117,  13'd626,  -13'd322,  -13'd542,  13'd329,  -13'd675,  13'd353,  
-13'd405,  13'd351,  -13'd333,  13'd637,  -13'd294,  -13'd105,  13'd306,  13'd52,  13'd508,  13'd157,  13'd422,  -13'd244,  13'd322,  -13'd843,  -13'd196,  -13'd122,  
13'd157,  13'd529,  13'd330,  -13'd179,  13'd27,  13'd281,  -13'd191,  -13'd750,  13'd414,  13'd421,  13'd179,  13'd546,  13'd183,  -13'd642,  -13'd38,  13'd157,  
13'd29,  13'd237,  13'd222,  13'd448,  -13'd260,  13'd114,  13'd43,  -13'd126,  13'd899,  13'd62,  13'd253,  -13'd669,  13'd442,  -13'd19,  13'd594,  13'd89,  
13'd754,  -13'd152,  -13'd262,  -13'd4,  -13'd225,  13'd100,  13'd596,  -13'd31,  -13'd291,  -13'd193,  13'd777,  -13'd298,  13'd447,  13'd538,  -13'd652,  -13'd509,  
13'd270,  13'd282,  -13'd536,  -13'd33,  13'd126,  -13'd69,  -13'd259,  -13'd18,  13'd314,  -13'd263,  13'd260,  -13'd46,  -13'd491,  -13'd42,  -13'd147,  -13'd354,  

-13'd261,  13'd869,  13'd686,  13'd208,  -13'd204,  13'd310,  13'd315,  -13'd892,  13'd405,  -13'd594,  -13'd881,  13'd381,  -13'd386,  13'd385,  -13'd343,  -13'd275,  
-13'd91,  -13'd54,  13'd1072,  -13'd972,  13'd115,  -13'd219,  -13'd98,  -13'd18,  13'd186,  -13'd181,  13'd190,  -13'd377,  13'd60,  13'd1167,  13'd45,  -13'd470,  
-13'd946,  13'd216,  13'd351,  -13'd69,  -13'd364,  13'd198,  -13'd239,  13'd35,  13'd73,  -13'd464,  13'd344,  13'd240,  -13'd829,  13'd1172,  -13'd153,  -13'd780,  
13'd178,  13'd10,  -13'd503,  13'd288,  -13'd130,  13'd599,  13'd240,  -13'd163,  13'd263,  13'd369,  -13'd705,  13'd239,  -13'd473,  13'd377,  -13'd500,  -13'd59,  
13'd574,  13'd294,  -13'd119,  13'd438,  -13'd243,  13'd122,  13'd489,  13'd24,  13'd673,  -13'd342,  -13'd78,  13'd362,  13'd585,  13'd568,  13'd42,  13'd520,  
13'd89,  13'd692,  13'd92,  13'd158,  -13'd622,  -13'd305,  13'd430,  13'd542,  -13'd383,  13'd933,  -13'd298,  13'd284,  -13'd344,  13'd932,  13'd561,  13'd241,  
13'd335,  13'd51,  13'd907,  -13'd563,  -13'd306,  -13'd795,  -13'd597,  13'd264,  13'd573,  -13'd79,  -13'd137,  -13'd387,  13'd534,  13'd1061,  13'd551,  13'd592,  
13'd69,  -13'd622,  13'd655,  -13'd24,  -13'd27,  -13'd45,  -13'd556,  13'd288,  13'd519,  13'd98,  13'd350,  -13'd338,  -13'd224,  13'd77,  -13'd670,  -13'd635,  
-13'd402,  13'd347,  13'd531,  -13'd240,  13'd125,  13'd569,  -13'd272,  13'd101,  -13'd64,  13'd412,  -13'd462,  13'd414,  -13'd331,  -13'd183,  13'd144,  13'd215,  
13'd580,  -13'd551,  -13'd403,  13'd48,  -13'd190,  13'd332,  -13'd161,  -13'd629,  13'd299,  -13'd1015,  -13'd255,  -13'd232,  -13'd642,  13'd193,  -13'd277,  13'd364,  
13'd814,  -13'd130,  -13'd19,  13'd828,  -13'd351,  13'd1244,  -13'd811,  13'd372,  13'd308,  13'd76,  13'd520,  -13'd229,  13'd1198,  13'd399,  -13'd125,  13'd347,  
-13'd220,  13'd708,  13'd120,  13'd347,  -13'd541,  13'd670,  -13'd144,  13'd865,  13'd295,  13'd562,  -13'd99,  -13'd123,  13'd255,  -13'd349,  13'd101,  -13'd728,  
13'd307,  -13'd80,  -13'd29,  13'd542,  -13'd141,  13'd813,  13'd300,  13'd277,  -13'd67,  -13'd209,  13'd850,  13'd31,  13'd779,  -13'd838,  -13'd421,  13'd22,  
-13'd56,  13'd136,  -13'd475,  13'd96,  13'd40,  -13'd467,  -13'd259,  -13'd461,  -13'd7,  -13'd581,  13'd792,  13'd420,  13'd31,  -13'd135,  13'd134,  -13'd156,  
-13'd247,  -13'd540,  -13'd90,  -13'd193,  -13'd219,  13'd49,  13'd362,  13'd314,  -13'd396,  -13'd471,  -13'd411,  -13'd37,  13'd1087,  -13'd129,  -13'd128,  13'd918,  
13'd233,  13'd791,  -13'd337,  13'd19,  13'd1485,  13'd301,  -13'd269,  -13'd379,  -13'd292,  13'd277,  -13'd117,  13'd853,  13'd412,  -13'd112,  13'd155,  13'd787,  
-13'd730,  -13'd107,  -13'd145,  -13'd24,  13'd351,  -13'd957,  13'd285,  13'd253,  -13'd149,  13'd160,  13'd165,  13'd162,  13'd211,  -13'd572,  -13'd287,  13'd202,  
-13'd113,  -13'd511,  13'd360,  13'd257,  13'd488,  -13'd291,  13'd288,  -13'd663,  13'd402,  13'd53,  -13'd208,  13'd160,  -13'd86,  13'd206,  -13'd553,  13'd53,  
13'd660,  13'd196,  13'd431,  13'd363,  -13'd327,  -13'd264,  13'd250,  -13'd59,  13'd520,  13'd742,  13'd601,  -13'd235,  -13'd65,  13'd625,  13'd48,  13'd726,  
-13'd360,  13'd408,  13'd254,  -13'd295,  -13'd483,  -13'd518,  -13'd758,  -13'd389,  -13'd779,  -13'd7,  -13'd196,  -13'd305,  -13'd498,  -13'd515,  13'd394,  13'd612,  
13'd295,  13'd729,  -13'd183,  -13'd465,  13'd472,  13'd251,  13'd155,  -13'd288,  13'd593,  -13'd668,  -13'd452,  13'd875,  -13'd630,  -13'd252,  -13'd268,  -13'd303,  
13'd170,  -13'd678,  -13'd122,  -13'd466,  13'd22,  -13'd245,  13'd842,  -13'd529,  -13'd61,  -13'd266,  -13'd166,  13'd66,  -13'd617,  -13'd230,  13'd603,  -13'd419,  
13'd655,  -13'd39,  13'd254,  -13'd246,  13'd318,  -13'd595,  13'd55,  -13'd228,  13'd72,  13'd262,  -13'd534,  -13'd485,  -13'd600,  13'd681,  -13'd156,  -13'd132,  
-13'd216,  13'd9,  -13'd53,  -13'd54,  -13'd363,  13'd57,  -13'd394,  13'd346,  13'd307,  13'd15,  -13'd44,  -13'd1,  -13'd408,  13'd948,  13'd608,  -13'd86,  
13'd129,  -13'd505,  13'd1163,  13'd659,  13'd94,  13'd59,  13'd320,  13'd446,  -13'd183,  -13'd461,  -13'd429,  13'd154,  13'd594,  -13'd266,  13'd1200,  13'd679,  

13'd302,  -13'd7,  -13'd497,  -13'd856,  -13'd837,  13'd764,  13'd620,  13'd147,  13'd800,  -13'd547,  13'd193,  13'd197,  -13'd133,  13'd463,  -13'd466,  -13'd43,  
-13'd96,  -13'd772,  -13'd481,  13'd232,  -13'd66,  13'd375,  -13'd475,  -13'd711,  -13'd125,  -13'd572,  13'd193,  -13'd18,  -13'd89,  -13'd274,  13'd600,  13'd354,  
13'd444,  13'd105,  -13'd351,  13'd368,  -13'd545,  13'd401,  -13'd247,  13'd221,  13'd164,  -13'd156,  13'd120,  -13'd515,  -13'd236,  -13'd587,  -13'd146,  -13'd24,  
-13'd599,  -13'd3,  -13'd69,  13'd573,  13'd408,  13'd264,  -13'd361,  -13'd455,  -13'd195,  13'd124,  13'd397,  -13'd224,  13'd431,  -13'd1477,  13'd204,  13'd370,  
-13'd901,  -13'd892,  13'd286,  13'd125,  13'd505,  -13'd603,  -13'd317,  13'd312,  -13'd178,  -13'd505,  13'd352,  -13'd290,  13'd390,  13'd541,  -13'd188,  13'd966,  
13'd208,  13'd357,  -13'd132,  13'd554,  -13'd35,  13'd292,  -13'd683,  -13'd279,  -13'd692,  13'd982,  -13'd796,  13'd7,  -13'd322,  -13'd270,  13'd18,  13'd252,  
13'd289,  -13'd112,  13'd195,  13'd809,  -13'd673,  -13'd25,  -13'd1155,  13'd504,  13'd541,  -13'd366,  -13'd163,  -13'd676,  13'd741,  13'd63,  13'd489,  13'd310,  
-13'd665,  13'd82,  13'd16,  -13'd396,  -13'd359,  13'd64,  13'd181,  13'd50,  13'd802,  13'd867,  13'd1344,  -13'd278,  13'd135,  -13'd81,  -13'd275,  -13'd14,  
-13'd1409,  -13'd657,  -13'd150,  -13'd387,  -13'd423,  -13'd259,  13'd406,  13'd477,  13'd147,  13'd1017,  13'd24,  -13'd117,  13'd139,  -13'd270,  13'd526,  13'd201,  
-13'd496,  13'd4,  13'd207,  -13'd214,  -13'd569,  13'd265,  -13'd358,  -13'd124,  13'd433,  13'd297,  13'd528,  13'd365,  13'd311,  -13'd838,  13'd110,  13'd342,  
13'd429,  13'd8,  -13'd430,  -13'd82,  13'd494,  -13'd184,  -13'd1602,  -13'd3,  13'd483,  13'd565,  13'd357,  -13'd277,  13'd385,  -13'd53,  -13'd110,  -13'd17,  
-13'd320,  13'd561,  13'd313,  -13'd531,  13'd35,  13'd232,  -13'd477,  13'd859,  13'd415,  13'd167,  -13'd422,  13'd436,  -13'd65,  13'd139,  -13'd107,  -13'd399,  
13'd402,  -13'd347,  -13'd610,  13'd218,  13'd691,  13'd244,  13'd116,  -13'd549,  -13'd51,  -13'd308,  13'd267,  13'd321,  13'd652,  -13'd370,  13'd350,  -13'd579,  
-13'd333,  13'd595,  13'd90,  -13'd329,  13'd245,  -13'd572,  -13'd84,  13'd264,  -13'd358,  13'd318,  13'd617,  -13'd107,  -13'd341,  -13'd84,  -13'd121,  -13'd201,  
13'd378,  13'd419,  -13'd213,  -13'd231,  13'd149,  13'd638,  13'd385,  13'd190,  13'd93,  -13'd14,  13'd255,  -13'd341,  13'd716,  -13'd272,  13'd241,  -13'd140,  
13'd321,  -13'd23,  13'd129,  13'd474,  13'd866,  13'd137,  13'd841,  -13'd400,  13'd957,  13'd614,  -13'd29,  -13'd222,  13'd212,  13'd457,  13'd363,  13'd731,  
13'd799,  13'd410,  13'd145,  13'd111,  -13'd222,  13'd132,  -13'd357,  -13'd169,  13'd207,  13'd364,  13'd373,  13'd915,  13'd1002,  13'd100,  13'd194,  13'd476,  
-13'd165,  -13'd2,  -13'd84,  13'd568,  13'd173,  -13'd453,  13'd89,  -13'd455,  13'd232,  13'd754,  -13'd202,  -13'd443,  -13'd1,  -13'd614,  -13'd313,  13'd229,  
-13'd226,  -13'd205,  -13'd471,  -13'd287,  13'd253,  -13'd417,  13'd57,  -13'd347,  -13'd83,  13'd2,  -13'd522,  -13'd336,  -13'd511,  -13'd347,  13'd427,  13'd539,  
13'd480,  -13'd674,  13'd728,  13'd349,  -13'd180,  13'd717,  13'd21,  -13'd222,  13'd280,  13'd1376,  13'd124,  -13'd586,  13'd131,  13'd547,  -13'd109,  13'd195,  
13'd77,  -13'd119,  -13'd136,  13'd526,  13'd275,  13'd362,  13'd587,  13'd807,  13'd616,  13'd491,  13'd384,  -13'd493,  13'd659,  -13'd224,  -13'd29,  -13'd246,  
13'd444,  -13'd966,  -13'd369,  -13'd493,  13'd471,  -13'd381,  -13'd269,  13'd111,  -13'd226,  -13'd165,  13'd49,  -13'd180,  13'd255,  13'd380,  -13'd49,  13'd108,  
-13'd617,  -13'd424,  -13'd433,  -13'd141,  13'd75,  13'd51,  -13'd335,  -13'd498,  13'd98,  13'd98,  -13'd252,  13'd848,  -13'd222,  13'd78,  13'd122,  -13'd88,  
13'd242,  -13'd137,  -13'd511,  13'd193,  13'd284,  -13'd171,  -13'd312,  -13'd29,  13'd419,  -13'd445,  13'd111,  -13'd333,  -13'd262,  13'd352,  -13'd311,  13'd465,  
-13'd26,  13'd85,  13'd111,  13'd387,  -13'd2,  13'd362,  -13'd37,  13'd408,  -13'd158,  -13'd243,  13'd425,  -13'd75,  13'd96,  -13'd309,  13'd420,  13'd714,  

-13'd445,  13'd243,  13'd488,  -13'd510,  13'd483,  -13'd820,  13'd192,  -13'd925,  13'd326,  13'd265,  13'd312,  -13'd452,  13'd265,  13'd923,  13'd195,  13'd581,  
-13'd689,  -13'd655,  13'd521,  -13'd42,  13'd66,  -13'd241,  13'd666,  -13'd708,  13'd49,  -13'd538,  13'd226,  13'd177,  -13'd366,  13'd963,  -13'd215,  13'd324,  
13'd552,  -13'd314,  13'd609,  -13'd447,  -13'd1157,  13'd64,  -13'd52,  -13'd247,  -13'd478,  -13'd315,  13'd705,  -13'd785,  -13'd581,  13'd1230,  13'd288,  -13'd407,  
13'd459,  13'd286,  -13'd490,  -13'd713,  -13'd336,  -13'd124,  13'd532,  13'd507,  13'd297,  -13'd136,  -13'd247,  13'd33,  13'd609,  -13'd608,  13'd460,  -13'd75,  
13'd261,  13'd1705,  -13'd960,  13'd615,  -13'd186,  13'd211,  13'd367,  -13'd64,  -13'd74,  13'd24,  13'd852,  13'd177,  13'd1159,  13'd249,  13'd36,  13'd1059,  
-13'd606,  -13'd186,  13'd377,  -13'd265,  -13'd618,  -13'd514,  13'd533,  -13'd307,  -13'd402,  -13'd180,  13'd752,  -13'd30,  13'd210,  13'd543,  13'd231,  13'd268,  
13'd344,  13'd25,  -13'd190,  13'd289,  13'd478,  -13'd511,  13'd804,  13'd340,  -13'd11,  -13'd38,  13'd793,  13'd230,  13'd30,  13'd393,  -13'd668,  -13'd612,  
13'd117,  -13'd729,  13'd270,  -13'd821,  13'd127,  13'd72,  -13'd248,  13'd34,  13'd1038,  -13'd28,  13'd150,  13'd129,  -13'd81,  -13'd307,  -13'd641,  -13'd372,  
13'd413,  13'd1004,  13'd49,  13'd283,  13'd108,  -13'd8,  -13'd396,  13'd1215,  13'd318,  13'd274,  13'd791,  -13'd124,  -13'd154,  -13'd291,  13'd187,  -13'd567,  
13'd87,  13'd196,  13'd254,  -13'd16,  13'd431,  13'd589,  -13'd58,  13'd712,  -13'd35,  13'd1217,  13'd214,  13'd95,  -13'd157,  13'd414,  13'd910,  13'd8,  
13'd645,  13'd55,  13'd329,  -13'd349,  -13'd1429,  13'd624,  13'd1053,  -13'd275,  -13'd676,  13'd303,  13'd330,  13'd385,  -13'd160,  -13'd81,  13'd346,  13'd845,  
-13'd243,  13'd347,  13'd476,  13'd72,  13'd315,  -13'd332,  13'd204,  13'd250,  13'd5,  13'd36,  -13'd409,  -13'd170,  -13'd184,  13'd827,  -13'd94,  -13'd156,  
-13'd462,  13'd197,  13'd39,  -13'd479,  13'd352,  -13'd443,  -13'd282,  -13'd173,  -13'd245,  -13'd281,  -13'd5,  -13'd101,  13'd457,  -13'd170,  -13'd505,  13'd211,  
-13'd391,  -13'd367,  -13'd773,  -13'd163,  13'd197,  -13'd304,  -13'd869,  -13'd553,  -13'd358,  13'd711,  -13'd377,  13'd158,  -13'd177,  -13'd749,  13'd489,  13'd652,  
-13'd194,  13'd82,  13'd374,  -13'd10,  13'd467,  -13'd154,  -13'd654,  -13'd342,  13'd247,  13'd127,  13'd286,  13'd307,  -13'd45,  -13'd281,  13'd943,  13'd393,  
13'd85,  13'd222,  13'd829,  13'd88,  -13'd361,  13'd226,  -13'd110,  13'd1125,  13'd104,  13'd31,  13'd195,  -13'd2,  -13'd27,  13'd41,  13'd383,  13'd129,  
-13'd249,  13'd379,  13'd203,  13'd820,  -13'd526,  13'd187,  -13'd61,  13'd6,  -13'd896,  -13'd427,  -13'd204,  -13'd698,  -13'd625,  13'd171,  13'd229,  -13'd760,  
13'd306,  -13'd542,  13'd323,  13'd275,  13'd576,  -13'd361,  13'd2,  13'd172,  13'd431,  -13'd594,  -13'd26,  -13'd98,  13'd529,  13'd517,  -13'd350,  -13'd646,  
13'd85,  -13'd144,  -13'd642,  -13'd183,  13'd790,  13'd573,  13'd69,  -13'd85,  13'd125,  13'd3,  13'd702,  13'd245,  13'd6,  13'd10,  -13'd61,  13'd27,  
13'd542,  13'd960,  13'd864,  -13'd551,  13'd175,  13'd124,  13'd375,  13'd72,  13'd146,  -13'd235,  -13'd33,  13'd510,  13'd178,  -13'd266,  13'd256,  -13'd5,  
-13'd858,  -13'd74,  -13'd79,  -13'd106,  -13'd228,  13'd446,  -13'd172,  13'd88,  13'd66,  -13'd39,  -13'd298,  13'd389,  -13'd455,  13'd235,  -13'd343,  13'd78,  
-13'd836,  -13'd306,  13'd181,  13'd518,  13'd389,  13'd860,  13'd733,  13'd41,  13'd533,  -13'd126,  13'd405,  -13'd133,  13'd695,  -13'd265,  -13'd119,  13'd45,  
-13'd494,  13'd110,  -13'd269,  13'd101,  13'd135,  13'd533,  13'd201,  13'd194,  13'd728,  -13'd188,  13'd790,  13'd120,  -13'd168,  -13'd337,  -13'd423,  13'd480,  
13'd942,  13'd103,  13'd877,  13'd176,  -13'd48,  -13'd257,  -13'd599,  13'd617,  -13'd78,  13'd250,  13'd485,  13'd491,  13'd282,  13'd158,  -13'd909,  -13'd438,  
13'd697,  13'd39,  13'd516,  -13'd73,  13'd340,  -13'd136,  13'd379,  -13'd237,  13'd777,  13'd342,  -13'd311,  13'd1149,  13'd374,  -13'd688,  13'd5,  -13'd127,  

-13'd815,  -13'd108,  -13'd417,  13'd79,  13'd267,  13'd85,  -13'd673,  13'd628,  -13'd421,  13'd138,  -13'd134,  -13'd700,  13'd1095,  -13'd149,  -13'd130,  -13'd712,  
-13'd253,  13'd373,  13'd63,  -13'd27,  13'd399,  13'd459,  -13'd379,  13'd18,  13'd254,  13'd224,  -13'd680,  -13'd130,  13'd362,  -13'd136,  13'd417,  13'd83,  
-13'd535,  -13'd141,  13'd858,  13'd113,  -13'd699,  13'd357,  13'd336,  -13'd585,  13'd49,  -13'd392,  13'd136,  -13'd393,  -13'd295,  13'd673,  13'd495,  13'd796,  
-13'd187,  -13'd374,  13'd44,  13'd909,  -13'd795,  -13'd581,  -13'd405,  -13'd11,  13'd894,  13'd219,  13'd544,  13'd20,  -13'd549,  13'd84,  13'd117,  -13'd234,  
-13'd19,  -13'd560,  13'd390,  -13'd270,  13'd733,  -13'd525,  -13'd438,  -13'd474,  -13'd158,  -13'd285,  13'd563,  13'd106,  -13'd174,  13'd106,  -13'd83,  13'd61,  
-13'd664,  -13'd202,  -13'd956,  13'd555,  13'd379,  -13'd778,  -13'd175,  -13'd798,  13'd120,  -13'd536,  13'd502,  -13'd235,  13'd240,  -13'd35,  -13'd638,  13'd308,  
-13'd439,  -13'd490,  -13'd843,  13'd478,  13'd993,  -13'd414,  -13'd403,  -13'd173,  -13'd285,  13'd373,  -13'd401,  13'd573,  13'd678,  -13'd398,  -13'd25,  13'd459,  
-13'd108,  13'd142,  13'd95,  13'd295,  13'd189,  -13'd206,  -13'd13,  -13'd76,  -13'd334,  13'd12,  13'd375,  13'd260,  13'd493,  -13'd112,  -13'd981,  -13'd51,  
-13'd50,  13'd60,  13'd210,  -13'd430,  -13'd229,  13'd487,  -13'd412,  -13'd401,  -13'd367,  13'd370,  13'd430,  13'd84,  13'd228,  13'd884,  -13'd22,  -13'd78,  
13'd278,  13'd855,  13'd666,  13'd438,  -13'd194,  -13'd543,  13'd509,  -13'd47,  13'd426,  13'd399,  13'd106,  13'd8,  -13'd504,  13'd523,  13'd880,  -13'd286,  
-13'd394,  13'd267,  -13'd617,  -13'd710,  -13'd458,  13'd572,  -13'd925,  13'd255,  13'd720,  -13'd435,  13'd806,  13'd226,  -13'd92,  -13'd40,  13'd434,  13'd434,  
13'd441,  13'd89,  13'd15,  13'd178,  13'd216,  13'd424,  -13'd367,  -13'd645,  13'd225,  13'd1121,  13'd103,  13'd112,  13'd271,  -13'd670,  -13'd598,  13'd951,  
13'd319,  13'd273,  -13'd782,  13'd261,  13'd925,  -13'd709,  13'd83,  13'd312,  -13'd337,  13'd333,  13'd648,  13'd612,  13'd66,  -13'd259,  13'd9,  13'd797,  
13'd135,  13'd386,  13'd372,  13'd174,  13'd399,  -13'd234,  13'd367,  13'd328,  13'd587,  13'd599,  13'd571,  -13'd266,  -13'd470,  13'd83,  -13'd684,  -13'd877,  
13'd502,  13'd219,  13'd86,  13'd416,  -13'd792,  13'd488,  13'd173,  -13'd138,  13'd229,  -13'd511,  -13'd598,  -13'd85,  13'd639,  -13'd447,  -13'd1008,  -13'd91,  
13'd36,  -13'd160,  -13'd493,  -13'd81,  -13'd750,  -13'd269,  -13'd524,  -13'd264,  13'd331,  -13'd32,  13'd751,  -13'd245,  -13'd156,  -13'd609,  13'd60,  13'd370,  
-13'd463,  13'd22,  -13'd663,  13'd318,  13'd275,  -13'd24,  -13'd484,  13'd744,  -13'd249,  13'd129,  13'd401,  13'd506,  13'd232,  -13'd348,  13'd214,  13'd505,  
13'd360,  13'd622,  -13'd733,  13'd212,  13'd365,  13'd151,  -13'd137,  13'd138,  13'd163,  -13'd468,  13'd407,  13'd526,  13'd295,  13'd418,  -13'd308,  -13'd136,  
13'd196,  -13'd220,  -13'd688,  13'd880,  13'd147,  -13'd396,  -13'd90,  13'd44,  13'd196,  -13'd407,  13'd788,  -13'd298,  13'd503,  -13'd14,  13'd106,  13'd466,  
13'd414,  -13'd345,  -13'd629,  13'd338,  13'd680,  13'd605,  -13'd120,  -13'd358,  13'd481,  -13'd67,  13'd77,  13'd43,  13'd1231,  13'd125,  -13'd59,  13'd121,  
-13'd79,  -13'd341,  -13'd173,  -13'd508,  -13'd147,  -13'd16,  13'd748,  -13'd724,  -13'd685,  13'd532,  13'd285,  -13'd294,  13'd438,  13'd18,  13'd360,  13'd430,  
-13'd51,  13'd767,  13'd287,  -13'd218,  13'd61,  -13'd912,  -13'd154,  -13'd2,  -13'd18,  -13'd257,  13'd685,  -13'd322,  13'd3,  -13'd1027,  13'd113,  13'd292,  
13'd421,  13'd281,  -13'd369,  -13'd36,  13'd517,  -13'd170,  -13'd254,  -13'd340,  -13'd410,  13'd1028,  -13'd364,  -13'd27,  13'd348,  -13'd190,  13'd385,  -13'd471,  
-13'd625,  13'd905,  -13'd86,  13'd324,  13'd31,  -13'd496,  -13'd239,  -13'd50,  -13'd50,  13'd76,  13'd56,  -13'd811,  13'd756,  13'd126,  -13'd260,  -13'd505,  
13'd94,  13'd670,  13'd229,  -13'd315,  -13'd114,  13'd451,  -13'd930,  13'd427,  13'd199,  13'd664,  -13'd672,  13'd251,  -13'd320,  -13'd326,  13'd119,  -13'd217,  

13'd214,  13'd3,  -13'd481,  -13'd54,  -13'd64,  13'd116,  13'd6,  -13'd233,  13'd518,  -13'd231,  -13'd301,  13'd277,  13'd408,  -13'd127,  -13'd558,  13'd316,  
13'd559,  -13'd221,  13'd250,  13'd317,  -13'd544,  13'd253,  -13'd62,  13'd46,  -13'd751,  13'd345,  -13'd603,  -13'd17,  -13'd605,  -13'd501,  -13'd687,  -13'd366,  
-13'd229,  -13'd471,  -13'd149,  -13'd48,  13'd64,  13'd81,  -13'd16,  -13'd374,  13'd256,  -13'd346,  -13'd108,  -13'd457,  -13'd279,  -13'd253,  -13'd276,  13'd252,  
-13'd426,  -13'd282,  -13'd365,  13'd1,  -13'd31,  -13'd104,  13'd131,  13'd247,  13'd196,  -13'd360,  -13'd143,  13'd308,  -13'd273,  -13'd656,  -13'd63,  -13'd283,  
13'd64,  13'd337,  13'd378,  -13'd371,  -13'd106,  -13'd370,  -13'd117,  13'd6,  13'd210,  13'd15,  -13'd599,  -13'd27,  13'd49,  13'd244,  13'd544,  13'd305,  
-13'd239,  -13'd262,  -13'd236,  -13'd324,  13'd78,  13'd268,  -13'd468,  -13'd423,  13'd12,  -13'd721,  13'd358,  13'd64,  -13'd355,  13'd352,  -13'd200,  -13'd184,  
13'd487,  13'd5,  13'd298,  -13'd391,  13'd333,  -13'd491,  -13'd35,  -13'd341,  -13'd273,  -13'd315,  13'd264,  13'd22,  13'd503,  -13'd138,  13'd157,  13'd271,  
13'd70,  -13'd435,  -13'd343,  -13'd192,  13'd240,  -13'd100,  -13'd847,  13'd406,  -13'd183,  13'd18,  13'd174,  -13'd654,  13'd505,  -13'd104,  -13'd115,  -13'd530,  
13'd600,  -13'd225,  13'd23,  -13'd20,  13'd85,  13'd663,  -13'd554,  13'd225,  -13'd487,  -13'd375,  -13'd193,  13'd148,  13'd434,  -13'd322,  13'd440,  13'd265,  
13'd514,  -13'd104,  13'd280,  13'd726,  -13'd70,  -13'd331,  -13'd712,  13'd583,  13'd81,  -13'd736,  -13'd186,  -13'd75,  -13'd107,  -13'd45,  13'd467,  13'd463,  
-13'd55,  13'd64,  -13'd135,  -13'd273,  -13'd720,  13'd146,  -13'd383,  -13'd183,  -13'd357,  -13'd765,  -13'd156,  13'd35,  13'd113,  -13'd84,  13'd403,  -13'd670,  
13'd499,  -13'd181,  13'd490,  13'd328,  -13'd851,  13'd356,  -13'd157,  13'd185,  -13'd716,  13'd657,  13'd346,  13'd36,  13'd310,  -13'd383,  13'd43,  13'd89,  
13'd7,  -13'd342,  -13'd563,  -13'd49,  13'd24,  -13'd738,  13'd120,  -13'd158,  13'd342,  13'd151,  -13'd259,  13'd182,  -13'd126,  13'd89,  13'd309,  13'd252,  
-13'd232,  13'd259,  -13'd378,  -13'd7,  -13'd28,  -13'd358,  -13'd328,  -13'd438,  -13'd735,  -13'd728,  -13'd354,  -13'd391,  -13'd409,  13'd119,  -13'd338,  -13'd135,  
-13'd476,  13'd34,  -13'd541,  -13'd373,  -13'd300,  -13'd109,  -13'd39,  -13'd695,  -13'd32,  -13'd322,  -13'd633,  -13'd161,  13'd14,  -13'd77,  13'd295,  13'd35,  
-13'd201,  -13'd13,  -13'd75,  -13'd50,  13'd159,  -13'd282,  -13'd260,  13'd87,  13'd439,  -13'd250,  -13'd355,  -13'd221,  -13'd316,  -13'd130,  13'd313,  13'd495,  
13'd334,  13'd615,  13'd271,  -13'd430,  -13'd90,  13'd474,  -13'd759,  -13'd20,  13'd130,  -13'd181,  13'd162,  13'd69,  -13'd44,  13'd205,  -13'd382,  13'd342,  
-13'd729,  13'd31,  -13'd77,  13'd79,  -13'd539,  13'd500,  13'd292,  -13'd13,  -13'd596,  -13'd435,  -13'd1,  -13'd281,  -13'd528,  -13'd247,  13'd181,  -13'd61,  
13'd530,  -13'd51,  -13'd334,  13'd376,  13'd530,  13'd290,  -13'd53,  -13'd365,  13'd472,  -13'd194,  -13'd290,  13'd61,  13'd674,  13'd124,  13'd206,  -13'd35,  
13'd598,  -13'd645,  -13'd265,  -13'd385,  -13'd193,  -13'd230,  -13'd343,  -13'd42,  -13'd413,  13'd355,  13'd89,  13'd74,  -13'd156,  13'd550,  -13'd276,  13'd356,  
-13'd148,  13'd248,  -13'd12,  13'd576,  -13'd743,  13'd307,  13'd191,  -13'd155,  13'd66,  -13'd600,  -13'd74,  -13'd486,  13'd283,  -13'd551,  -13'd601,  -13'd737,  
-13'd209,  13'd46,  -13'd317,  13'd597,  13'd186,  -13'd766,  -13'd112,  -13'd342,  13'd192,  13'd380,  13'd221,  13'd245,  -13'd844,  -13'd222,  -13'd271,  -13'd501,  
-13'd143,  13'd25,  -13'd605,  -13'd323,  13'd110,  13'd149,  -13'd392,  -13'd367,  13'd63,  -13'd605,  13'd573,  -13'd718,  -13'd238,  -13'd612,  13'd404,  -13'd532,  
-13'd372,  -13'd243,  13'd134,  -13'd176,  -13'd383,  13'd706,  -13'd53,  -13'd234,  -13'd131,  13'd456,  -13'd359,  13'd326,  -13'd464,  -13'd172,  13'd150,  -13'd431,  
13'd97,  13'd169,  13'd26,  -13'd115,  13'd176,  -13'd410,  13'd4,  -13'd454,  13'd645,  -13'd386,  13'd515,  -13'd349,  -13'd644,  -13'd78,  13'd54,  -13'd255,  

-13'd443,  -13'd64,  -13'd308,  -13'd10,  13'd181,  13'd432,  13'd166,  -13'd474,  -13'd818,  13'd2,  -13'd151,  13'd422,  -13'd249,  -13'd413,  -13'd532,  -13'd356,  
13'd56,  -13'd169,  -13'd739,  -13'd45,  -13'd248,  13'd150,  -13'd142,  13'd211,  -13'd33,  13'd155,  13'd192,  13'd370,  -13'd507,  -13'd998,  -13'd222,  13'd158,  
-13'd856,  -13'd414,  -13'd261,  -13'd194,  13'd1043,  13'd263,  -13'd400,  -13'd493,  -13'd637,  13'd321,  13'd140,  -13'd40,  13'd822,  -13'd1616,  -13'd133,  -13'd13,  
-13'd974,  -13'd835,  13'd327,  13'd236,  13'd56,  -13'd794,  -13'd73,  13'd131,  -13'd504,  -13'd10,  -13'd213,  13'd370,  13'd118,  -13'd18,  13'd188,  -13'd280,  
-13'd184,  -13'd232,  -13'd86,  -13'd444,  13'd717,  -13'd288,  -13'd325,  13'd547,  13'd357,  -13'd294,  13'd139,  13'd288,  -13'd310,  -13'd189,  -13'd195,  -13'd83,  
-13'd735,  13'd307,  13'd42,  -13'd423,  -13'd541,  -13'd713,  -13'd3,  13'd376,  13'd695,  -13'd320,  13'd957,  13'd335,  13'd239,  13'd217,  13'd107,  13'd134,  
13'd91,  13'd486,  13'd411,  13'd68,  13'd86,  -13'd614,  13'd296,  -13'd486,  -13'd27,  13'd589,  -13'd715,  13'd422,  13'd449,  -13'd431,  13'd719,  13'd435,  
-13'd425,  -13'd441,  -13'd725,  -13'd15,  13'd338,  -13'd271,  13'd76,  -13'd383,  -13'd194,  -13'd176,  13'd99,  13'd642,  13'd533,  -13'd1100,  13'd559,  -13'd13,  
13'd252,  -13'd184,  -13'd207,  13'd176,  -13'd171,  -13'd79,  13'd412,  13'd388,  13'd483,  13'd71,  13'd85,  13'd250,  13'd555,  13'd495,  13'd297,  13'd785,  
13'd463,  13'd339,  13'd205,  13'd857,  13'd46,  13'd369,  13'd85,  13'd264,  -13'd357,  -13'd920,  -13'd45,  -13'd22,  13'd161,  13'd306,  -13'd339,  -13'd12,  
13'd117,  13'd51,  -13'd445,  -13'd180,  13'd271,  -13'd114,  -13'd973,  13'd49,  13'd363,  13'd285,  -13'd765,  -13'd347,  13'd737,  13'd375,  13'd334,  13'd268,  
-13'd22,  13'd297,  -13'd437,  13'd130,  -13'd86,  -13'd417,  -13'd734,  -13'd164,  -13'd598,  13'd235,  13'd641,  -13'd587,  -13'd50,  13'd444,  13'd323,  -13'd34,  
13'd544,  -13'd686,  13'd205,  13'd586,  -13'd443,  13'd294,  -13'd503,  -13'd28,  -13'd609,  13'd230,  13'd253,  13'd770,  -13'd118,  -13'd1252,  13'd38,  -13'd222,  
13'd413,  -13'd918,  -13'd189,  -13'd75,  13'd695,  -13'd366,  13'd289,  -13'd405,  13'd21,  13'd675,  -13'd340,  13'd181,  13'd330,  13'd98,  13'd92,  13'd484,  
-13'd291,  -13'd425,  -13'd182,  -13'd537,  13'd571,  -13'd92,  13'd462,  -13'd943,  -13'd345,  13'd300,  13'd291,  -13'd536,  -13'd38,  -13'd29,  13'd118,  13'd926,  
-13'd813,  -13'd263,  -13'd805,  -13'd292,  13'd530,  -13'd728,  -13'd633,  -13'd333,  -13'd107,  -13'd80,  -13'd295,  -13'd222,  -13'd454,  -13'd462,  -13'd407,  13'd273,  
13'd611,  13'd269,  -13'd148,  13'd636,  13'd1045,  -13'd409,  -13'd546,  -13'd594,  13'd626,  13'd364,  -13'd490,  13'd72,  13'd69,  -13'd929,  -13'd253,  13'd146,  
-13'd192,  13'd383,  13'd384,  13'd406,  -13'd617,  13'd459,  -13'd205,  13'd518,  13'd118,  -13'd188,  13'd158,  -13'd103,  -13'd276,  -13'd1307,  13'd513,  -13'd120,  
13'd189,  13'd470,  -13'd219,  -13'd159,  -13'd92,  -13'd188,  13'd260,  13'd229,  13'd850,  -13'd346,  -13'd29,  13'd274,  13'd231,  13'd562,  -13'd233,  -13'd253,  
-13'd54,  13'd84,  -13'd193,  -13'd141,  -13'd855,  -13'd459,  13'd533,  -13'd872,  13'd566,  -13'd260,  13'd264,  -13'd830,  -13'd457,  -13'd362,  -13'd497,  -13'd369,  
13'd241,  -13'd104,  -13'd342,  -13'd722,  -13'd352,  -13'd102,  13'd397,  -13'd357,  13'd955,  -13'd45,  13'd774,  13'd447,  13'd496,  -13'd782,  13'd358,  13'd53,  
13'd839,  -13'd518,  -13'd197,  -13'd37,  13'd241,  13'd121,  -13'd102,  13'd248,  13'd490,  13'd378,  13'd216,  13'd492,  -13'd200,  -13'd101,  -13'd498,  -13'd56,  
13'd155,  13'd377,  13'd544,  -13'd42,  -13'd768,  -13'd59,  13'd447,  13'd545,  13'd774,  13'd893,  13'd268,  13'd391,  13'd584,  13'd360,  13'd96,  -13'd219,  
13'd197,  -13'd254,  13'd400,  -13'd122,  -13'd389,  -13'd382,  13'd233,  -13'd70,  -13'd266,  -13'd456,  13'd125,  13'd485,  13'd233,  13'd801,  -13'd528,  13'd510,  
-13'd33,  -13'd474,  13'd460,  -13'd257,  -13'd645,  13'd93,  13'd154,  -13'd67,  13'd675,  -13'd222,  13'd3,  -13'd171,  -13'd77,  13'd254,  -13'd107,  -13'd374,  

13'd494,  -13'd471,  -13'd119,  -13'd836,  -13'd159,  -13'd149,  -13'd599,  13'd11,  13'd416,  13'd517,  -13'd43,  -13'd186,  -13'd44,  13'd6,  13'd214,  13'd69,  
13'd615,  -13'd136,  13'd185,  -13'd319,  13'd514,  13'd85,  -13'd347,  -13'd442,  13'd399,  -13'd845,  -13'd202,  -13'd630,  -13'd660,  -13'd138,  -13'd147,  13'd355,  
-13'd483,  -13'd238,  -13'd105,  13'd591,  -13'd265,  13'd358,  13'd566,  13'd621,  -13'd834,  -13'd575,  -13'd344,  -13'd354,  -13'd591,  13'd347,  13'd56,  13'd206,  
13'd129,  13'd421,  13'd226,  -13'd236,  13'd195,  -13'd55,  13'd573,  -13'd270,  -13'd295,  13'd75,  13'd262,  -13'd145,  13'd616,  -13'd286,  13'd95,  -13'd265,  
-13'd132,  13'd460,  13'd190,  -13'd495,  -13'd535,  13'd541,  -13'd148,  -13'd52,  -13'd377,  13'd176,  13'd61,  -13'd588,  13'd88,  -13'd50,  -13'd561,  13'd433,  
-13'd204,  13'd8,  -13'd300,  -13'd198,  -13'd331,  -13'd537,  -13'd536,  -13'd163,  13'd248,  -13'd479,  -13'd529,  -13'd19,  13'd594,  -13'd314,  -13'd409,  -13'd391,  
13'd195,  -13'd354,  13'd709,  13'd577,  -13'd225,  -13'd97,  -13'd402,  -13'd648,  13'd493,  -13'd0,  -13'd295,  13'd130,  13'd21,  13'd55,  -13'd650,  -13'd847,  
-13'd139,  13'd323,  13'd176,  13'd95,  13'd261,  -13'd145,  -13'd360,  -13'd218,  -13'd575,  -13'd106,  -13'd90,  13'd392,  13'd568,  13'd181,  -13'd404,  -13'd220,  
13'd369,  -13'd318,  -13'd219,  -13'd359,  13'd701,  13'd550,  -13'd353,  -13'd557,  -13'd385,  -13'd694,  13'd350,  -13'd356,  13'd48,  13'd171,  -13'd362,  -13'd146,  
-13'd400,  -13'd382,  13'd469,  -13'd483,  13'd398,  -13'd148,  13'd523,  -13'd484,  13'd187,  -13'd49,  -13'd108,  -13'd336,  -13'd618,  13'd260,  -13'd460,  13'd291,  
-13'd460,  -13'd509,  13'd170,  13'd294,  13'd56,  -13'd114,  -13'd164,  -13'd182,  -13'd90,  -13'd454,  -13'd893,  -13'd533,  13'd311,  13'd460,  13'd333,  -13'd78,  
13'd300,  13'd455,  -13'd329,  -13'd264,  -13'd184,  13'd23,  13'd416,  -13'd137,  -13'd118,  -13'd583,  13'd154,  13'd225,  13'd192,  -13'd395,  -13'd783,  13'd14,  
13'd115,  -13'd604,  13'd4,  -13'd317,  -13'd149,  -13'd349,  13'd224,  -13'd449,  13'd157,  13'd40,  -13'd20,  -13'd153,  -13'd471,  -13'd140,  -13'd151,  13'd609,  
-13'd369,  -13'd657,  13'd68,  -13'd45,  13'd260,  -13'd390,  -13'd85,  -13'd489,  -13'd749,  -13'd225,  -13'd408,  13'd100,  -13'd598,  -13'd131,  13'd14,  13'd189,  
-13'd232,  -13'd269,  -13'd35,  -13'd194,  13'd105,  13'd9,  13'd379,  13'd15,  13'd647,  -13'd23,  13'd232,  -13'd379,  -13'd18,  13'd164,  13'd637,  -13'd187,  
13'd217,  13'd414,  13'd376,  13'd305,  -13'd583,  13'd489,  13'd726,  -13'd265,  13'd510,  -13'd184,  -13'd264,  -13'd308,  13'd273,  -13'd719,  13'd12,  -13'd702,  
13'd238,  -13'd21,  -13'd435,  13'd136,  -13'd161,  -13'd365,  13'd71,  13'd551,  -13'd54,  13'd416,  13'd591,  -13'd652,  13'd384,  -13'd628,  13'd385,  13'd298,  
-13'd117,  -13'd563,  -13'd834,  13'd505,  13'd143,  -13'd242,  13'd322,  -13'd554,  13'd365,  13'd301,  -13'd161,  13'd106,  -13'd375,  13'd117,  -13'd220,  -13'd21,  
-13'd743,  -13'd208,  -13'd112,  13'd44,  13'd12,  -13'd303,  -13'd234,  13'd39,  -13'd137,  -13'd162,  13'd173,  13'd666,  -13'd543,  -13'd33,  13'd5,  13'd26,  
-13'd724,  13'd284,  13'd588,  -13'd399,  -13'd435,  13'd26,  -13'd542,  13'd441,  -13'd688,  13'd28,  13'd395,  -13'd110,  13'd155,  -13'd127,  13'd265,  -13'd340,  
-13'd52,  -13'd705,  -13'd506,  -13'd7,  -13'd208,  -13'd300,  -13'd429,  -13'd683,  13'd283,  -13'd116,  -13'd56,  -13'd270,  -13'd603,  13'd358,  -13'd222,  -13'd41,  
13'd210,  13'd549,  13'd99,  -13'd39,  13'd222,  -13'd76,  13'd98,  -13'd176,  13'd658,  -13'd11,  13'd364,  13'd255,  -13'd4,  13'd253,  13'd109,  -13'd0,  
13'd445,  -13'd206,  -13'd54,  -13'd770,  13'd142,  -13'd220,  13'd436,  -13'd225,  13'd20,  13'd208,  -13'd542,  -13'd277,  -13'd8,  13'd121,  -13'd179,  -13'd697,  
13'd156,  -13'd78,  13'd237,  -13'd305,  13'd28,  -13'd418,  13'd650,  -13'd375,  -13'd184,  -13'd8,  13'd168,  -13'd129,  -13'd467,  -13'd193,  -13'd348,  -13'd237,  
13'd552,  13'd147,  13'd244,  -13'd117,  -13'd312,  13'd275,  13'd383,  13'd100,  13'd110,  -13'd454,  13'd426,  -13'd183,  13'd126,  -13'd202,  -13'd494,  -13'd359,  

13'd118,  -13'd318,  13'd332,  -13'd299,  -13'd489,  -13'd80,  -13'd385,  -13'd124,  -13'd319,  13'd526,  13'd317,  -13'd14,  13'd396,  -13'd159,  -13'd384,  -13'd774,  
-13'd208,  13'd319,  -13'd463,  -13'd448,  -13'd600,  13'd374,  13'd329,  -13'd744,  13'd18,  -13'd447,  -13'd191,  -13'd298,  13'd49,  -13'd82,  13'd106,  13'd210,  
-13'd19,  13'd726,  13'd140,  -13'd221,  -13'd4,  13'd392,  13'd83,  -13'd409,  13'd543,  13'd607,  13'd8,  -13'd256,  -13'd650,  -13'd273,  -13'd407,  13'd44,  
13'd138,  -13'd635,  -13'd556,  13'd560,  13'd435,  13'd627,  13'd329,  -13'd530,  -13'd232,  13'd312,  -13'd589,  13'd252,  -13'd302,  -13'd753,  -13'd685,  -13'd263,  
13'd395,  -13'd121,  -13'd135,  -13'd467,  13'd574,  13'd183,  13'd62,  -13'd237,  13'd199,  13'd323,  -13'd116,  -13'd129,  -13'd644,  -13'd20,  13'd373,  13'd168,  
-13'd514,  13'd553,  -13'd699,  -13'd676,  -13'd921,  13'd36,  -13'd34,  -13'd635,  13'd307,  -13'd664,  -13'd642,  -13'd354,  -13'd397,  13'd175,  -13'd142,  -13'd140,  
-13'd515,  -13'd262,  -13'd502,  13'd402,  -13'd162,  -13'd727,  -13'd561,  -13'd307,  -13'd278,  -13'd926,  -13'd499,  -13'd519,  -13'd422,  -13'd275,  -13'd194,  -13'd465,  
-13'd329,  -13'd7,  -13'd661,  -13'd424,  -13'd193,  -13'd310,  13'd445,  -13'd352,  -13'd597,  13'd677,  -13'd406,  -13'd255,  13'd36,  -13'd875,  -13'd471,  13'd273,  
-13'd31,  -13'd405,  13'd89,  -13'd602,  -13'd536,  -13'd430,  -13'd24,  -13'd494,  13'd262,  -13'd147,  -13'd346,  13'd45,  13'd37,  -13'd449,  13'd56,  -13'd79,  
13'd5,  -13'd809,  13'd457,  -13'd305,  13'd367,  13'd297,  13'd512,  -13'd116,  13'd69,  13'd265,  -13'd315,  -13'd25,  13'd213,  -13'd127,  13'd474,  13'd85,  
-13'd677,  13'd316,  -13'd125,  -13'd585,  -13'd315,  -13'd416,  -13'd430,  13'd345,  13'd245,  13'd500,  -13'd326,  -13'd466,  -13'd90,  13'd137,  13'd517,  -13'd134,  
-13'd385,  -13'd250,  -13'd614,  -13'd113,  -13'd5,  13'd144,  -13'd256,  -13'd948,  13'd292,  -13'd214,  -13'd248,  13'd192,  -13'd272,  -13'd495,  13'd3,  -13'd97,  
13'd149,  -13'd677,  -13'd334,  13'd251,  13'd357,  13'd120,  13'd145,  -13'd132,  -13'd841,  -13'd346,  13'd155,  -13'd64,  -13'd307,  13'd114,  -13'd331,  13'd65,  
13'd131,  -13'd176,  -13'd943,  13'd21,  13'd201,  -13'd169,  13'd20,  13'd84,  -13'd79,  13'd177,  13'd142,  -13'd228,  -13'd312,  13'd516,  13'd71,  13'd98,  
-13'd223,  -13'd81,  -13'd168,  -13'd161,  13'd217,  -13'd312,  -13'd91,  -13'd471,  13'd30,  -13'd494,  -13'd669,  13'd335,  13'd434,  13'd246,  -13'd394,  13'd84,  
-13'd569,  13'd121,  -13'd14,  -13'd558,  13'd4,  -13'd165,  13'd22,  -13'd560,  -13'd239,  -13'd208,  -13'd57,  -13'd375,  -13'd210,  13'd147,  -13'd189,  13'd275,  
-13'd1,  -13'd14,  -13'd19,  -13'd160,  13'd39,  -13'd608,  -13'd53,  13'd113,  -13'd672,  13'd402,  13'd21,  -13'd667,  -13'd619,  13'd375,  13'd607,  13'd261,  
-13'd647,  -13'd311,  13'd213,  -13'd197,  -13'd143,  -13'd562,  -13'd177,  13'd462,  13'd793,  13'd260,  -13'd793,  -13'd435,  -13'd310,  13'd77,  13'd121,  -13'd313,  
-13'd402,  13'd473,  -13'd992,  -13'd337,  -13'd324,  -13'd116,  13'd45,  -13'd209,  -13'd618,  -13'd387,  -13'd680,  13'd197,  -13'd34,  -13'd243,  -13'd585,  -13'd105,  
13'd89,  -13'd666,  -13'd206,  -13'd568,  -13'd41,  -13'd315,  -13'd266,  -13'd609,  -13'd103,  -13'd148,  -13'd420,  -13'd701,  13'd100,  -13'd23,  13'd159,  13'd345,  
-13'd412,  -13'd16,  -13'd343,  -13'd910,  -13'd205,  -13'd169,  13'd178,  13'd205,  13'd208,  -13'd761,  -13'd113,  -13'd202,  13'd121,  -13'd16,  13'd84,  -13'd225,  
13'd425,  -13'd225,  -13'd429,  -13'd482,  -13'd276,  13'd357,  13'd280,  -13'd649,  13'd334,  13'd98,  13'd190,  13'd33,  13'd80,  13'd239,  13'd8,  -13'd495,  
13'd227,  -13'd226,  -13'd661,  13'd406,  13'd345,  13'd297,  13'd116,  -13'd415,  -13'd210,  13'd108,  13'd590,  13'd43,  -13'd41,  -13'd548,  13'd0,  13'd320,  
13'd384,  -13'd497,  -13'd318,  -13'd186,  -13'd327,  -13'd516,  -13'd338,  -13'd268,  13'd337,  -13'd502,  -13'd132,  -13'd5,  -13'd30,  13'd22,  13'd53,  13'd119,  
-13'd149,  13'd282,  -13'd144,  -13'd183,  13'd245,  -13'd356,  -13'd632,  -13'd411,  13'd91,  -13'd694,  13'd522,  -13'd292,  -13'd624,  -13'd293,  13'd199,  13'd256,  

13'd394,  13'd505,  13'd1117,  13'd668,  -13'd95,  13'd49,  -13'd736,  13'd46,  -13'd189,  13'd412,  -13'd198,  -13'd72,  13'd482,  13'd365,  13'd644,  -13'd372,  
13'd531,  13'd313,  -13'd326,  -13'd20,  13'd734,  -13'd702,  13'd296,  -13'd290,  13'd1143,  -13'd537,  -13'd84,  13'd832,  13'd216,  -13'd501,  -13'd503,  13'd93,  
13'd383,  13'd715,  -13'd540,  -13'd2,  -13'd397,  13'd749,  13'd162,  -13'd352,  -13'd553,  -13'd228,  -13'd368,  13'd11,  13'd130,  13'd912,  13'd100,  13'd381,  
13'd55,  13'd34,  13'd520,  -13'd30,  13'd135,  -13'd779,  -13'd105,  -13'd272,  13'd271,  -13'd98,  -13'd67,  13'd293,  13'd272,  13'd861,  -13'd435,  13'd375,  
13'd130,  13'd811,  -13'd844,  -13'd257,  13'd107,  -13'd117,  13'd536,  -13'd248,  13'd508,  13'd504,  13'd386,  13'd560,  -13'd202,  13'd849,  13'd154,  13'd14,  
-13'd389,  -13'd284,  13'd663,  -13'd85,  13'd158,  13'd46,  13'd508,  13'd676,  -13'd174,  13'd630,  13'd542,  -13'd130,  13'd289,  13'd315,  -13'd168,  13'd68,  
-13'd527,  -13'd271,  13'd504,  -13'd176,  -13'd580,  13'd137,  13'd383,  13'd151,  -13'd57,  13'd390,  13'd79,  -13'd111,  13'd311,  -13'd341,  13'd3,  -13'd717,  
13'd71,  13'd599,  -13'd39,  -13'd419,  13'd111,  -13'd435,  13'd296,  -13'd587,  13'd73,  -13'd1,  -13'd376,  13'd789,  13'd705,  -13'd158,  13'd67,  -13'd110,  
13'd422,  13'd364,  -13'd401,  13'd221,  13'd137,  -13'd27,  13'd137,  -13'd1015,  13'd72,  -13'd1051,  -13'd483,  13'd278,  -13'd42,  13'd529,  -13'd385,  13'd265,  
-13'd57,  13'd332,  -13'd1025,  -13'd380,  13'd625,  -13'd352,  13'd405,  -13'd373,  13'd373,  -13'd171,  13'd407,  13'd399,  13'd626,  -13'd296,  13'd47,  -13'd196,  
13'd254,  13'd23,  13'd183,  13'd528,  -13'd534,  -13'd120,  13'd523,  13'd64,  -13'd16,  13'd416,  13'd362,  -13'd117,  13'd91,  13'd323,  13'd721,  13'd496,  
13'd217,  13'd12,  13'd220,  -13'd208,  -13'd60,  -13'd78,  13'd556,  13'd415,  13'd419,  13'd284,  13'd692,  -13'd251,  13'd83,  -13'd740,  13'd96,  -13'd221,  
13'd698,  -13'd758,  13'd431,  13'd922,  13'd401,  13'd513,  -13'd795,  13'd228,  13'd60,  13'd482,  13'd115,  13'd511,  13'd450,  13'd700,  13'd524,  13'd399,  
13'd598,  -13'd976,  -13'd511,  -13'd380,  13'd570,  -13'd194,  13'd332,  -13'd534,  -13'd399,  -13'd191,  -13'd516,  13'd329,  13'd567,  13'd206,  -13'd125,  -13'd430,  
13'd171,  -13'd638,  -13'd417,  13'd56,  -13'd298,  13'd2,  -13'd444,  -13'd606,  13'd5,  13'd528,  -13'd362,  13'd309,  -13'd243,  13'd524,  -13'd88,  13'd667,  
13'd236,  -13'd38,  13'd256,  -13'd355,  13'd596,  -13'd745,  13'd854,  -13'd53,  -13'd390,  13'd27,  13'd61,  13'd297,  13'd307,  13'd20,  -13'd32,  13'd575,  
13'd370,  -13'd502,  -13'd607,  -13'd2,  -13'd435,  13'd118,  13'd350,  13'd170,  13'd713,  13'd639,  -13'd448,  -13'd373,  -13'd252,  13'd649,  -13'd101,  13'd235,  
-13'd346,  13'd463,  -13'd278,  13'd350,  -13'd387,  13'd254,  13'd175,  -13'd127,  -13'd31,  -13'd440,  13'd587,  13'd494,  13'd197,  -13'd550,  -13'd296,  13'd68,  
-13'd86,  -13'd451,  -13'd205,  13'd242,  13'd851,  -13'd86,  -13'd51,  -13'd5,  -13'd124,  -13'd184,  13'd559,  -13'd373,  -13'd116,  -13'd184,  -13'd81,  -13'd530,  
-13'd171,  -13'd471,  -13'd470,  13'd322,  13'd935,  13'd82,  13'd205,  13'd154,  13'd209,  13'd654,  13'd14,  13'd554,  13'd148,  -13'd391,  -13'd204,  13'd612,  
13'd421,  13'd782,  -13'd240,  -13'd705,  -13'd118,  -13'd421,  -13'd13,  -13'd264,  -13'd891,  -13'd549,  13'd64,  -13'd30,  -13'd114,  13'd479,  13'd0,  -13'd551,  
-13'd338,  -13'd313,  13'd901,  13'd52,  -13'd216,  -13'd476,  -13'd660,  13'd394,  -13'd798,  -13'd721,  -13'd752,  -13'd294,  -13'd338,  13'd1538,  -13'd302,  -13'd197,  
-13'd305,  13'd374,  13'd225,  -13'd113,  13'd170,  13'd1,  -13'd0,  -13'd85,  -13'd353,  -13'd515,  -13'd42,  -13'd222,  -13'd112,  13'd626,  13'd604,  -13'd560,  
-13'd539,  -13'd436,  -13'd608,  -13'd459,  -13'd409,  13'd734,  -13'd248,  13'd166,  -13'd259,  -13'd465,  13'd393,  13'd116,  13'd331,  13'd854,  13'd1001,  13'd804,  
-13'd1111,  13'd485,  13'd77,  13'd672,  -13'd153,  -13'd213,  13'd41,  -13'd66,  -13'd760,  -13'd107,  13'd558,  13'd315,  -13'd345,  -13'd103,  13'd988,  13'd315
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule



module bias_fc2_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC2-1][0:`OUTPUT_NUM_FC2-1][`WD_BIAS:0] weight	 = {
		24'd376858,  24'd432250,  24'd29999,  -24'd21180,  24'd203900,  -24'd35257,  24'd214653,  -24'd285062,  24'd149942,  24'd172424,  24'd241287,  24'd324760,  24'd306054,  24'd109385,  24'd386902,  24'd1789,  
24'd28800,  24'd347429,  24'd509845,  24'd403218,  24'd55283,  24'd293083,  -24'd21746,  -24'd254371,  -24'd400996,  -24'd132702,  -24'd107502,  -24'd140243,  -24'd206663,  -24'd140441,  24'd143746,  24'd39439,  
24'd236044,  24'd268803,  24'd150150,  24'd385287,  -24'd213047,  24'd26023,  -24'd343539,  24'd332436,  -24'd397889,  -24'd209506,  -24'd133163,  24'd243649,  -24'd9532,  24'd307082,  -24'd132963,  -24'd159572,  
-24'd53911,  24'd55608,  -24'd63297,  24'd287278,  24'd231376,  24'd227915,  -24'd149391,  24'd406123,  -24'd279679,  24'd37076,  24'd251134,  24'd110896,  -24'd132970,  24'd307661,  24'd327144,  24'd66815,  
24'd131364,  24'd119973,  -24'd302322,  24'd158931,  24'd47008,  -24'd154135,  -24'd42487,  24'd329397,  24'd366838,  24'd373655,  24'd391455,  24'd142308,  24'd61661,  24'd27682,  24'd173948,  -24'd11642,  
24'd233626,  -24'd79977,  24'd87200,  24'd305044
	 };
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule


module wieght_fc2_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2*`OUTPUT_BATCH_FC2)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC1*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC2*`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2-1][0:`OUTPUT_NUM_FC2-1][0:`OUTPUT_NUM_FC1-1][`WD:0] weight	 = {
13'd84,  -13'd337,  -13'd547,  13'd779,  13'd1037,  -13'd210,  13'd435,  13'd816,  -13'd690,  -13'd128,  -13'd783,  13'd810,  -13'd559,  -13'd188,  13'd935,  13'd291,  
13'd434,  -13'd59,  -13'd39,  13'd467,  13'd511,  -13'd953,  13'd62,  13'd967,  13'd42,  -13'd98,  -13'd235,  -13'd92,  -13'd342,  13'd283,  13'd208,  -13'd429,  
13'd381,  13'd663,  -13'd519,  13'd298,  -13'd185,  13'd167,  13'd259,  13'd713,  -13'd179,  -13'd723,  13'd200,  13'd343,  13'd598,  13'd162,  -13'd860,  -13'd328,  
-13'd200,  13'd191,  13'd153,  13'd383,  -13'd377,  13'd268,  -13'd615,  13'd48,  13'd496,  -13'd513,  13'd32,  -13'd301,  13'd68,  13'd689,  -13'd173,  13'd464,  
13'd52,  13'd541,  13'd338,  -13'd399,  -13'd122,  -13'd451,  -13'd221,  13'd112,  13'd348,  13'd882,  -13'd436,  -13'd584,  13'd372,  -13'd184,  -13'd536,  13'd447,  
-13'd126,  -13'd78,  13'd222,  13'd33,  13'd317,  -13'd671,  -13'd495,  13'd129,  -13'd586,  13'd273,  -13'd697,  -13'd642,  13'd377,  13'd258,  13'd675,  -13'd330,  
-13'd48,  -13'd423,  -13'd148,  13'd1219,  -13'd161,  -13'd476,  13'd61,  -13'd127,  -13'd581,  -13'd311,  -13'd760,  13'd853,  -13'd493,  -13'd476,  13'd219,  13'd434,  
13'd370,  13'd159,  -13'd598,  -13'd29,  13'd384,  -13'd79,  -13'd717,  -13'd471,  
-13'd361,  -13'd460,  13'd148,  13'd46,  -13'd72,  -13'd401,  -13'd724,  -13'd822,  13'd135,  13'd113,  13'd188,  -13'd899,  13'd8,  13'd149,  13'd682,  13'd415,  
-13'd27,  -13'd258,  13'd678,  -13'd294,  -13'd53,  13'd693,  13'd158,  -13'd333,  13'd151,  -13'd621,  -13'd203,  -13'd340,  13'd364,  13'd432,  13'd409,  13'd20,  
-13'd213,  -13'd82,  13'd846,  13'd362,  13'd203,  13'd135,  -13'd151,  -13'd48,  13'd552,  -13'd756,  13'd291,  13'd144,  13'd337,  -13'd20,  -13'd495,  -13'd790,  
13'd185,  -13'd719,  -13'd65,  13'd212,  13'd795,  13'd450,  -13'd693,  -13'd286,  -13'd316,  13'd472,  -13'd410,  13'd437,  13'd673,  13'd286,  13'd157,  13'd137,  
13'd248,  13'd71,  13'd176,  13'd25,  -13'd443,  13'd82,  -13'd505,  13'd34,  -13'd678,  -13'd401,  13'd76,  -13'd129,  -13'd362,  -13'd526,  13'd207,  -13'd267,  
13'd36,  -13'd72,  13'd629,  -13'd187,  -13'd35,  -13'd498,  -13'd34,  13'd23,  -13'd15,  -13'd73,  -13'd502,  13'd460,  13'd591,  13'd434,  -13'd567,  13'd206,  
13'd653,  13'd619,  -13'd378,  13'd90,  13'd377,  -13'd197,  13'd370,  -13'd1114,  13'd546,  13'd88,  -13'd413,  -13'd747,  -13'd59,  13'd350,  -13'd694,  13'd602,  
13'd107,  -13'd45,  -13'd338,  -13'd21,  13'd502,  13'd145,  13'd704,  -13'd224,  
-13'd655,  -13'd323,  13'd328,  13'd474,  -13'd107,  13'd421,  13'd105,  13'd253,  -13'd470,  13'd14,  13'd37,  -13'd256,  13'd83,  13'd382,  -13'd35,  13'd383,  
-13'd481,  13'd196,  -13'd415,  13'd70,  13'd159,  13'd410,  -13'd129,  13'd239,  -13'd564,  -13'd538,  -13'd274,  13'd350,  -13'd117,  13'd218,  -13'd156,  13'd643,  
-13'd259,  13'd577,  13'd500,  13'd536,  -13'd536,  13'd687,  -13'd164,  13'd433,  13'd715,  13'd287,  -13'd275,  -13'd233,  -13'd192,  13'd803,  13'd149,  -13'd468,  
13'd66,  -13'd707,  13'd789,  13'd120,  13'd92,  -13'd983,  13'd609,  13'd262,  -13'd45,  13'd487,  13'd566,  13'd527,  13'd445,  -13'd241,  -13'd611,  -13'd143,  
-13'd400,  13'd79,  -13'd86,  -13'd284,  -13'd20,  -13'd339,  -13'd99,  13'd418,  -13'd127,  13'd320,  13'd523,  -13'd386,  -13'd699,  -13'd313,  13'd194,  -13'd583,  
13'd305,  -13'd631,  -13'd737,  -13'd185,  13'd443,  13'd198,  13'd534,  13'd283,  13'd41,  -13'd425,  13'd195,  -13'd370,  -13'd755,  13'd860,  13'd317,  -13'd25,  
-13'd574,  -13'd26,  13'd18,  -13'd40,  -13'd319,  13'd315,  -13'd558,  13'd597,  13'd57,  13'd445,  13'd248,  13'd186,  -13'd162,  -13'd25,  13'd529,  13'd280,  
13'd98,  13'd43,  13'd61,  -13'd101,  13'd961,  -13'd364,  -13'd31,  13'd338,  
13'd286,  -13'd74,  13'd183,  -13'd30,  13'd466,  13'd192,  13'd190,  -13'd495,  -13'd711,  13'd36,  -13'd740,  -13'd521,  13'd327,  13'd127,  13'd168,  13'd254,  
13'd658,  13'd304,  -13'd209,  -13'd609,  13'd305,  13'd343,  13'd570,  13'd92,  13'd395,  -13'd654,  13'd26,  -13'd1075,  13'd219,  13'd7,  13'd546,  13'd1031,  
13'd130,  13'd12,  13'd162,  13'd122,  13'd726,  -13'd271,  -13'd814,  13'd449,  -13'd288,  13'd193,  13'd351,  -13'd858,  13'd510,  13'd257,  -13'd1094,  -13'd302,  
-13'd195,  13'd654,  13'd733,  13'd63,  -13'd189,  13'd114,  13'd38,  -13'd24,  13'd415,  13'd582,  -13'd20,  13'd18,  13'd231,  -13'd358,  13'd168,  -13'd660,  
-13'd206,  13'd98,  -13'd215,  13'd653,  -13'd816,  13'd61,  -13'd933,  -13'd17,  13'd406,  -13'd704,  -13'd91,  13'd372,  -13'd772,  -13'd277,  13'd593,  13'd189,  
-13'd242,  -13'd363,  13'd406,  -13'd130,  -13'd540,  13'd221,  13'd153,  -13'd486,  -13'd247,  -13'd196,  13'd538,  -13'd333,  13'd258,  -13'd27,  13'd636,  -13'd151,  
13'd546,  -13'd60,  13'd139,  -13'd267,  13'd660,  13'd909,  -13'd131,  -13'd1710,  13'd116,  -13'd281,  -13'd368,  -13'd243,  13'd56,  -13'd1114,  -13'd516,  13'd705,  
13'd49,  13'd47,  13'd70,  -13'd703,  -13'd794,  -13'd350,  13'd139,  13'd731,  
-13'd391,  -13'd75,  -13'd528,  -13'd303,  13'd375,  13'd499,  13'd382,  -13'd189,  -13'd180,  13'd396,  -13'd767,  13'd416,  13'd385,  13'd302,  13'd153,  13'd26,  
13'd288,  -13'd75,  13'd397,  -13'd414,  -13'd43,  13'd516,  13'd297,  13'd41,  13'd256,  -13'd615,  -13'd94,  13'd454,  13'd158,  -13'd257,  13'd368,  -13'd289,  
-13'd448,  13'd455,  -13'd240,  -13'd77,  -13'd69,  13'd19,  -13'd161,  13'd823,  -13'd821,  -13'd63,  -13'd1185,  -13'd272,  13'd218,  13'd400,  13'd831,  13'd483,  
13'd445,  -13'd615,  -13'd666,  13'd651,  13'd94,  13'd597,  13'd245,  -13'd364,  -13'd189,  -13'd101,  13'd340,  -13'd202,  -13'd34,  13'd527,  13'd324,  -13'd331,  
13'd670,  -13'd273,  13'd372,  -13'd699,  13'd968,  -13'd169,  -13'd254,  13'd602,  13'd21,  -13'd2,  -13'd395,  -13'd6,  13'd161,  13'd69,  -13'd225,  13'd573,  
-13'd26,  -13'd383,  13'd589,  -13'd621,  -13'd205,  -13'd172,  -13'd149,  13'd77,  -13'd635,  13'd329,  13'd252,  13'd245,  13'd436,  -13'd525,  -13'd175,  -13'd126,  
-13'd233,  13'd138,  13'd317,  -13'd841,  -13'd22,  13'd2,  13'd443,  -13'd352,  -13'd133,  -13'd31,  -13'd330,  13'd1385,  13'd378,  -13'd220,  -13'd737,  -13'd146,  
13'd770,  -13'd338,  13'd617,  -13'd393,  -13'd198,  13'd434,  13'd34,  -13'd388,  
-13'd722,  -13'd33,  13'd666,  13'd52,  -13'd804,  13'd811,  13'd278,  -13'd613,  -13'd145,  13'd407,  13'd1101,  -13'd619,  -13'd388,  13'd4,  -13'd188,  -13'd75,  
-13'd77,  -13'd38,  -13'd369,  13'd297,  13'd169,  13'd448,  13'd593,  -13'd14,  -13'd57,  13'd101,  13'd452,  -13'd21,  -13'd333,  13'd582,  -13'd502,  -13'd85,  
-13'd409,  13'd195,  13'd97,  -13'd174,  13'd437,  13'd213,  -13'd476,  -13'd750,  13'd359,  13'd80,  -13'd237,  13'd703,  -13'd754,  13'd21,  -13'd148,  13'd224,  
13'd526,  13'd131,  13'd375,  13'd639,  13'd798,  13'd132,  13'd873,  13'd101,  -13'd1059,  13'd153,  -13'd400,  -13'd106,  13'd640,  13'd100,  13'd462,  -13'd594,  
-13'd215,  -13'd600,  -13'd545,  13'd265,  -13'd759,  13'd484,  -13'd44,  -13'd54,  13'd137,  13'd556,  13'd222,  13'd313,  -13'd571,  13'd104,  -13'd194,  13'd310,  
13'd351,  -13'd190,  13'd154,  -13'd828,  13'd295,  13'd834,  13'd252,  -13'd428,  -13'd69,  13'd31,  13'd452,  13'd75,  -13'd59,  13'd329,  13'd182,  13'd421,  
13'd506,  13'd287,  13'd493,  -13'd195,  13'd464,  -13'd477,  13'd687,  13'd490,  13'd82,  -13'd335,  13'd96,  -13'd215,  -13'd495,  13'd7,  13'd611,  -13'd259,  
-13'd23,  13'd571,  13'd1090,  13'd564,  -13'd212,  -13'd569,  -13'd438,  -13'd159,  
13'd242,  -13'd350,  13'd398,  -13'd309,  -13'd523,  -13'd680,  -13'd900,  13'd369,  -13'd937,  -13'd263,  -13'd666,  -13'd471,  -13'd335,  13'd415,  -13'd610,  13'd276,  
-13'd179,  13'd134,  13'd21,  -13'd189,  13'd354,  -13'd606,  -13'd93,  13'd370,  13'd413,  13'd455,  13'd409,  -13'd387,  -13'd134,  13'd94,  -13'd173,  13'd646,  
-13'd241,  13'd333,  13'd637,  13'd179,  13'd948,  -13'd259,  -13'd813,  -13'd670,  13'd2,  -13'd354,  -13'd152,  -13'd61,  -13'd638,  -13'd220,  -13'd544,  -13'd1588,  
13'd166,  13'd148,  -13'd22,  13'd391,  13'd117,  13'd300,  13'd334,  13'd408,  13'd441,  13'd269,  13'd171,  13'd661,  13'd567,  -13'd1199,  -13'd228,  13'd139,  
13'd125,  13'd136,  -13'd548,  -13'd407,  -13'd841,  13'd787,  -13'd101,  13'd120,  -13'd478,  13'd38,  13'd83,  -13'd380,  13'd408,  13'd412,  13'd276,  13'd110,  
-13'd240,  -13'd687,  -13'd64,  13'd343,  -13'd315,  -13'd601,  -13'd392,  -13'd183,  -13'd267,  13'd367,  13'd32,  -13'd406,  13'd267,  13'd578,  -13'd617,  13'd836,  
-13'd290,  -13'd449,  -13'd234,  -13'd282,  -13'd285,  13'd95,  13'd804,  13'd200,  -13'd520,  -13'd630,  -13'd20,  13'd328,  -13'd267,  -13'd356,  -13'd246,  13'd224,  
-13'd242,  13'd354,  -13'd808,  -13'd198,  13'd590,  13'd251,  13'd25,  -13'd221,  
13'd431,  -13'd127,  -13'd403,  -13'd475,  13'd478,  13'd263,  -13'd570,  -13'd142,  -13'd248,  -13'd262,  -13'd670,  13'd362,  13'd460,  -13'd91,  13'd715,  13'd104,  
13'd245,  13'd283,  -13'd236,  13'd42,  -13'd600,  13'd296,  -13'd238,  13'd957,  13'd231,  13'd834,  -13'd275,  -13'd627,  13'd734,  -13'd98,  13'd337,  13'd251,  
13'd310,  -13'd65,  -13'd196,  13'd94,  13'd695,  -13'd133,  13'd517,  -13'd51,  -13'd385,  -13'd288,  13'd56,  -13'd591,  13'd756,  13'd323,  -13'd138,  -13'd671,  
13'd124,  13'd343,  13'd337,  -13'd866,  -13'd90,  13'd241,  13'd728,  13'd179,  13'd43,  13'd422,  -13'd465,  13'd361,  13'd291,  13'd375,  13'd214,  -13'd336,  
13'd13,  13'd430,  13'd483,  -13'd152,  13'd202,  -13'd932,  13'd752,  13'd176,  13'd1042,  -13'd657,  -13'd85,  -13'd954,  13'd223,  -13'd245,  13'd157,  13'd308,  
-13'd80,  -13'd556,  -13'd741,  13'd583,  -13'd303,  -13'd74,  13'd128,  -13'd94,  -13'd905,  -13'd628,  13'd687,  13'd123,  13'd808,  -13'd672,  -13'd74,  -13'd361,  
-13'd296,  13'd403,  -13'd350,  13'd715,  13'd188,  -13'd428,  -13'd586,  -13'd186,  -13'd399,  13'd250,  -13'd158,  13'd157,  -13'd489,  -13'd190,  -13'd71,  13'd558,  
-13'd523,  -13'd308,  -13'd23,  13'd435,  13'd276,  13'd582,  -13'd29,  13'd417,  
13'd131,  13'd339,  -13'd455,  -13'd76,  -13'd541,  13'd261,  -13'd725,  -13'd47,  -13'd327,  -13'd483,  -13'd355,  13'd485,  -13'd154,  13'd966,  -13'd93,  13'd100,  
13'd134,  -13'd944,  13'd459,  13'd605,  13'd218,  13'd659,  13'd26,  -13'd393,  13'd31,  -13'd472,  -13'd332,  13'd35,  -13'd247,  13'd283,  -13'd913,  -13'd154,  
-13'd81,  13'd345,  -13'd284,  -13'd197,  13'd47,  13'd380,  -13'd764,  13'd206,  -13'd475,  13'd280,  -13'd433,  -13'd313,  13'd314,  13'd547,  -13'd354,  13'd199,  
13'd165,  13'd364,  -13'd187,  13'd115,  13'd594,  13'd316,  -13'd526,  13'd53,  -13'd336,  13'd437,  13'd698,  13'd158,  -13'd781,  13'd408,  13'd729,  13'd677,  
13'd390,  -13'd421,  13'd194,  -13'd438,  13'd402,  13'd139,  13'd88,  -13'd531,  13'd530,  13'd567,  -13'd299,  13'd102,  -13'd330,  -13'd340,  13'd178,  -13'd213,  
13'd328,  -13'd507,  13'd244,  -13'd53,  -13'd505,  -13'd104,  -13'd322,  13'd95,  -13'd218,  -13'd321,  -13'd60,  13'd142,  13'd281,  -13'd134,  -13'd299,  -13'd539,  
13'd79,  -13'd151,  13'd995,  -13'd428,  13'd169,  -13'd776,  -13'd74,  -13'd215,  13'd468,  -13'd307,  -13'd791,  13'd157,  -13'd270,  -13'd103,  -13'd133,  13'd457,  
13'd488,  13'd337,  13'd460,  13'd251,  -13'd684,  -13'd286,  13'd322,  13'd823,  
-13'd506,  13'd74,  -13'd243,  13'd121,  13'd388,  13'd89,  13'd352,  13'd1188,  -13'd390,  13'd206,  13'd488,  -13'd129,  -13'd180,  -13'd301,  13'd325,  -13'd176,  
-13'd155,  13'd503,  13'd393,  -13'd414,  13'd137,  -13'd285,  13'd384,  -13'd159,  13'd237,  13'd370,  -13'd81,  13'd235,  13'd75,  13'd653,  13'd286,  -13'd296,  
-13'd293,  13'd824,  -13'd434,  13'd271,  -13'd26,  -13'd1290,  -13'd455,  13'd616,  -13'd966,  -13'd326,  13'd247,  13'd836,  13'd1388,  13'd613,  -13'd64,  -13'd256,  
13'd621,  13'd192,  13'd681,  -13'd590,  13'd42,  -13'd408,  -13'd1897,  -13'd326,  13'd474,  13'd321,  -13'd111,  13'd1020,  13'd87,  -13'd228,  -13'd244,  13'd1075,  
13'd290,  -13'd117,  -13'd333,  -13'd373,  -13'd638,  13'd202,  -13'd245,  13'd378,  -13'd463,  -13'd116,  13'd498,  -13'd197,  13'd420,  -13'd123,  -13'd51,  -13'd309,  
-13'd606,  13'd953,  13'd69,  -13'd270,  -13'd149,  13'd594,  -13'd210,  -13'd228,  -13'd476,  13'd344,  -13'd84,  13'd50,  13'd523,  -13'd95,  13'd18,  13'd105,  
13'd138,  -13'd105,  -13'd541,  -13'd174,  13'd98,  -13'd1279,  13'd47,  -13'd658,  13'd155,  -13'd342,  -13'd161,  13'd52,  13'd291,  -13'd2,  -13'd429,  13'd833,  
-13'd543,  13'd620,  -13'd458,  13'd103,  13'd723,  13'd337,  -13'd100,  13'd340,  
-13'd396,  13'd818,  -13'd458,  13'd287,  13'd537,  13'd531,  -13'd331,  -13'd219,  -13'd168,  13'd185,  -13'd1913,  -13'd237,  13'd576,  13'd119,  13'd677,  13'd934,  
-13'd26,  -13'd161,  -13'd1219,  -13'd617,  13'd263,  13'd168,  13'd373,  13'd643,  13'd320,  -13'd811,  -13'd918,  -13'd687,  13'd533,  13'd86,  13'd1043,  13'd290,  
13'd172,  13'd584,  13'd752,  13'd622,  -13'd613,  13'd250,  13'd121,  13'd131,  -13'd31,  -13'd418,  13'd714,  -13'd203,  -13'd296,  13'd185,  13'd316,  -13'd1119,  
-13'd176,  -13'd600,  -13'd573,  13'd65,  -13'd54,  13'd721,  -13'd603,  13'd775,  13'd438,  13'd679,  -13'd1255,  13'd598,  -13'd266,  13'd488,  13'd311,  13'd3,  
13'd298,  -13'd189,  13'd581,  13'd108,  13'd8,  -13'd490,  13'd6,  13'd580,  -13'd264,  -13'd201,  -13'd412,  -13'd342,  13'd148,  13'd624,  -13'd720,  -13'd321,  
13'd341,  -13'd46,  13'd481,  -13'd57,  -13'd1244,  -13'd68,  -13'd276,  13'd365,  -13'd612,  -13'd295,  13'd56,  13'd464,  13'd744,  -13'd556,  -13'd731,  -13'd91,  
-13'd38,  -13'd621,  -13'd443,  -13'd146,  -13'd395,  13'd1085,  -13'd12,  -13'd710,  -13'd404,  13'd704,  13'd640,  13'd676,  13'd317,  -13'd826,  -13'd360,  13'd116,  
-13'd506,  -13'd307,  13'd210,  -13'd443,  -13'd159,  -13'd47,  13'd343,  13'd604,  
13'd135,  13'd287,  -13'd628,  13'd118,  13'd809,  13'd722,  -13'd167,  -13'd126,  -13'd49,  13'd960,  13'd321,  13'd532,  -13'd10,  13'd195,  -13'd125,  13'd1056,  
13'd611,  -13'd305,  -13'd150,  -13'd186,  -13'd63,  -13'd247,  13'd773,  13'd611,  13'd51,  13'd951,  -13'd277,  13'd376,  -13'd323,  13'd475,  13'd460,  -13'd679,  
-13'd445,  -13'd479,  13'd36,  13'd228,  -13'd72,  13'd553,  13'd238,  13'd186,  -13'd876,  13'd387,  -13'd102,  13'd368,  13'd826,  13'd123,  -13'd368,  13'd43,  
-13'd111,  -13'd64,  -13'd359,  13'd798,  13'd770,  13'd1041,  13'd631,  13'd760,  -13'd644,  -13'd413,  13'd28,  13'd491,  13'd648,  -13'd121,  13'd367,  13'd87,  
13'd1529,  -13'd151,  -13'd179,  -13'd278,  13'd207,  -13'd363,  13'd711,  13'd528,  13'd1079,  13'd553,  -13'd770,  13'd245,  -13'd536,  -13'd910,  -13'd240,  13'd39,  
-13'd106,  -13'd584,  -13'd808,  -13'd91,  -13'd62,  13'd449,  13'd85,  13'd108,  -13'd397,  -13'd356,  13'd748,  13'd151,  13'd289,  -13'd927,  -13'd166,  13'd99,  
-13'd77,  -13'd320,  13'd460,  13'd996,  -13'd849,  13'd1205,  13'd173,  -13'd226,  13'd233,  13'd481,  13'd643,  13'd311,  -13'd93,  13'd187,  13'd50,  13'd205,  
13'd510,  -13'd100,  13'd124,  -13'd695,  13'd246,  -13'd447,  -13'd325,  -13'd13,  
13'd224,  13'd100,  13'd77,  -13'd65,  13'd292,  13'd365,  -13'd99,  -13'd592,  -13'd417,  13'd217,  -13'd835,  13'd18,  13'd580,  13'd245,  -13'd294,  13'd245,  
13'd394,  13'd804,  -13'd442,  -13'd211,  13'd48,  -13'd367,  13'd664,  -13'd394,  -13'd132,  -13'd1101,  13'd9,  -13'd10,  13'd610,  13'd213,  -13'd232,  -13'd72,  
-13'd372,  13'd216,  13'd817,  -13'd262,  -13'd1042,  13'd805,  -13'd144,  -13'd701,  13'd263,  -13'd496,  -13'd836,  13'd316,  -13'd249,  13'd36,  13'd695,  13'd566,  
-13'd59,  -13'd1267,  13'd633,  -13'd298,  13'd198,  -13'd861,  -13'd40,  -13'd311,  13'd826,  -13'd58,  13'd538,  -13'd42,  -13'd308,  -13'd576,  -13'd468,  -13'd211,  
13'd696,  13'd269,  13'd583,  13'd838,  -13'd392,  -13'd429,  -13'd759,  13'd397,  -13'd579,  13'd656,  13'd363,  13'd568,  13'd562,  13'd703,  -13'd223,  13'd147,  
13'd36,  -13'd287,  -13'd472,  -13'd180,  13'd566,  13'd518,  13'd603,  13'd120,  13'd293,  -13'd42,  13'd658,  13'd459,  -13'd85,  13'd12,  13'd807,  13'd851,  
-13'd421,  13'd151,  13'd351,  13'd480,  -13'd305,  13'd479,  13'd223,  13'd541,  13'd289,  13'd233,  13'd689,  -13'd179,  -13'd248,  -13'd342,  13'd527,  -13'd424,  
13'd107,  -13'd399,  13'd359,  13'd660,  13'd215,  -13'd92,  -13'd631,  13'd54,  
13'd1258,  -13'd289,  13'd134,  13'd142,  13'd1048,  -13'd547,  -13'd941,  -13'd1075,  -13'd10,  -13'd101,  -13'd319,  -13'd584,  13'd321,  13'd337,  13'd193,  13'd445,  
13'd1155,  13'd694,  -13'd199,  -13'd85,  -13'd413,  13'd453,  13'd522,  13'd1140,  13'd329,  -13'd175,  -13'd408,  -13'd822,  -13'd483,  13'd347,  13'd25,  13'd9,  
13'd885,  -13'd21,  -13'd312,  13'd520,  13'd809,  13'd1175,  13'd320,  -13'd571,  13'd159,  13'd459,  -13'd36,  -13'd249,  -13'd193,  -13'd168,  13'd300,  -13'd1124,  
13'd8,  13'd288,  -13'd600,  13'd345,  13'd663,  -13'd112,  13'd427,  13'd831,  13'd203,  -13'd56,  -13'd35,  13'd433,  13'd556,  -13'd159,  -13'd484,  -13'd203,  
13'd455,  13'd261,  -13'd384,  13'd52,  -13'd376,  13'd360,  -13'd458,  -13'd712,  13'd369,  -13'd803,  13'd533,  -13'd873,  -13'd156,  13'd69,  -13'd324,  13'd566,  
13'd609,  -13'd4,  -13'd156,  13'd743,  13'd72,  13'd5,  -13'd75,  13'd841,  -13'd167,  13'd86,  13'd620,  -13'd381,  -13'd352,  13'd301,  -13'd414,  13'd161,  
13'd398,  13'd202,  -13'd232,  -13'd777,  -13'd438,  13'd376,  13'd495,  13'd595,  -13'd406,  13'd237,  13'd594,  -13'd833,  13'd597,  13'd755,  -13'd349,  13'd641,  
-13'd688,  -13'd177,  -13'd388,  -13'd30,  -13'd88,  -13'd112,  13'd325,  13'd194,  
13'd98,  -13'd223,  13'd581,  -13'd178,  13'd266,  -13'd200,  13'd349,  -13'd856,  -13'd402,  13'd235,  -13'd742,  -13'd527,  13'd593,  13'd77,  13'd1083,  -13'd141,  
13'd580,  13'd398,  -13'd734,  13'd167,  13'd41,  -13'd305,  13'd206,  13'd779,  13'd310,  -13'd127,  13'd142,  -13'd911,  13'd169,  -13'd617,  13'd368,  13'd1089,  
13'd514,  -13'd93,  13'd165,  13'd158,  13'd562,  13'd470,  13'd422,  -13'd224,  13'd64,  -13'd468,  -13'd55,  -13'd184,  13'd556,  -13'd683,  -13'd506,  -13'd981,  
-13'd355,  -13'd533,  -13'd445,  13'd1078,  -13'd164,  13'd608,  -13'd631,  13'd289,  13'd11,  13'd101,  -13'd586,  13'd738,  -13'd327,  -13'd364,  13'd375,  -13'd405,  
-13'd124,  13'd139,  13'd757,  13'd624,  -13'd173,  -13'd557,  13'd430,  13'd129,  -13'd457,  -13'd304,  -13'd490,  13'd127,  13'd230,  -13'd576,  13'd577,  -13'd267,  
13'd6,  -13'd109,  -13'd432,  13'd416,  13'd11,  -13'd629,  13'd557,  13'd240,  -13'd483,  13'd380,  13'd336,  -13'd180,  13'd632,  13'd91,  13'd194,  -13'd294,  
13'd280,  -13'd180,  -13'd564,  -13'd217,  -13'd376,  13'd1108,  13'd340,  13'd15,  -13'd163,  13'd207,  13'd460,  -13'd12,  13'd99,  -13'd599,  -13'd419,  13'd1175,  
13'd325,  -13'd268,  -13'd755,  13'd723,  13'd857,  -13'd41,  13'd527,  -13'd175,  
13'd32,  13'd181,  -13'd546,  -13'd212,  -13'd54,  -13'd186,  -13'd60,  -13'd142,  13'd771,  -13'd868,  -13'd7,  -13'd44,  13'd398,  13'd462,  -13'd20,  13'd583,  
13'd53,  -13'd142,  13'd696,  13'd144,  -13'd515,  -13'd102,  -13'd799,  13'd234,  -13'd484,  -13'd621,  -13'd163,  -13'd386,  -13'd347,  13'd292,  -13'd431,  -13'd222,  
13'd415,  13'd347,  13'd155,  -13'd262,  -13'd671,  13'd504,  -13'd486,  -13'd3,  -13'd253,  13'd713,  13'd32,  13'd201,  13'd6,  -13'd197,  -13'd360,  13'd53,  
-13'd42,  13'd15,  13'd255,  -13'd200,  13'd449,  13'd191,  -13'd86,  13'd290,  -13'd255,  13'd42,  -13'd266,  13'd223,  -13'd483,  -13'd363,  -13'd170,  -13'd47,  
-13'd641,  -13'd273,  13'd432,  13'd49,  -13'd576,  -13'd415,  13'd478,  13'd392,  13'd139,  -13'd241,  -13'd292,  13'd468,  13'd3,  -13'd207,  -13'd538,  13'd222,  
13'd774,  13'd351,  -13'd12,  -13'd280,  13'd533,  -13'd421,  13'd158,  13'd463,  13'd98,  13'd386,  13'd54,  -13'd285,  -13'd261,  -13'd42,  13'd379,  -13'd283,  
13'd478,  -13'd654,  13'd298,  13'd108,  -13'd374,  13'd191,  -13'd374,  -13'd310,  -13'd254,  -13'd164,  -13'd213,  -13'd470,  -13'd492,  -13'd218,  13'd148,  13'd134,  
-13'd96,  13'd197,  13'd256,  13'd115,  13'd81,  -13'd230,  -13'd312,  -13'd549,  
-13'd559,  -13'd152,  13'd182,  -13'd168,  -13'd125,  13'd67,  13'd312,  13'd268,  13'd148,  -13'd122,  13'd208,  13'd316,  -13'd443,  -13'd288,  13'd484,  -13'd135,  
-13'd536,  13'd473,  13'd303,  13'd391,  13'd229,  13'd219,  13'd164,  -13'd83,  -13'd324,  13'd272,  13'd91,  -13'd370,  -13'd606,  13'd413,  13'd288,  13'd399,  
-13'd63,  13'd269,  13'd90,  -13'd78,  13'd863,  -13'd199,  -13'd207,  -13'd275,  13'd770,  -13'd562,  13'd272,  13'd251,  13'd542,  13'd406,  13'd371,  13'd549,  
13'd158,  -13'd53,  13'd408,  -13'd332,  13'd106,  13'd927,  -13'd457,  13'd397,  -13'd644,  -13'd104,  -13'd198,  -13'd335,  13'd164,  13'd779,  13'd282,  13'd331,  
-13'd59,  13'd12,  -13'd131,  13'd194,  13'd302,  13'd593,  13'd665,  13'd292,  13'd79,  -13'd630,  13'd233,  -13'd67,  13'd59,  13'd245,  13'd49,  13'd636,  
13'd545,  13'd646,  -13'd141,  13'd791,  13'd395,  -13'd399,  13'd19,  -13'd753,  -13'd177,  -13'd580,  -13'd332,  13'd108,  13'd625,  -13'd486,  13'd58,  -13'd256,  
13'd788,  13'd307,  -13'd410,  -13'd389,  -13'd423,  -13'd785,  13'd181,  -13'd19,  -13'd305,  -13'd365,  -13'd283,  -13'd730,  -13'd138,  13'd220,  -13'd682,  13'd190,  
13'd46,  -13'd73,  13'd256,  13'd251,  -13'd509,  13'd68,  13'd2,  13'd538,  
-13'd568,  13'd360,  13'd36,  -13'd41,  13'd835,  -13'd323,  -13'd72,  -13'd1317,  13'd286,  13'd230,  13'd139,  -13'd164,  -13'd212,  -13'd428,  -13'd683,  -13'd666,  
13'd32,  13'd390,  -13'd171,  13'd653,  13'd110,  13'd480,  -13'd774,  13'd469,  13'd213,  13'd160,  13'd980,  13'd167,  13'd305,  13'd158,  13'd302,  -13'd691,  
-13'd233,  -13'd206,  -13'd94,  -13'd405,  -13'd654,  13'd400,  13'd491,  -13'd418,  13'd757,  -13'd105,  -13'd77,  13'd368,  -13'd72,  13'd204,  13'd796,  13'd402,  
13'd28,  13'd60,  -13'd566,  -13'd50,  13'd957,  13'd616,  -13'd993,  13'd199,  -13'd14,  13'd342,  13'd245,  -13'd476,  -13'd10,  13'd668,  13'd47,  -13'd183,  
-13'd188,  -13'd113,  -13'd150,  -13'd348,  13'd230,  13'd278,  13'd94,  -13'd468,  13'd61,  -13'd275,  -13'd129,  13'd122,  13'd776,  -13'd444,  -13'd164,  -13'd44,  
-13'd73,  13'd746,  13'd28,  13'd780,  -13'd486,  -13'd279,  -13'd444,  -13'd109,  13'd253,  13'd449,  13'd556,  -13'd336,  -13'd518,  13'd229,  13'd72,  -13'd450,  
13'd297,  -13'd305,  -13'd739,  13'd275,  -13'd145,  -13'd359,  13'd126,  -13'd1489,  -13'd305,  13'd513,  13'd482,  13'd722,  13'd523,  -13'd1057,  13'd127,  13'd152,  
13'd216,  -13'd139,  -13'd334,  -13'd391,  13'd102,  -13'd395,  -13'd340,  -13'd584,  
-13'd401,  -13'd36,  13'd659,  -13'd631,  13'd166,  -13'd225,  13'd128,  -13'd413,  13'd201,  13'd609,  13'd503,  -13'd233,  -13'd57,  -13'd17,  13'd327,  13'd550,  
-13'd247,  13'd49,  13'd782,  13'd102,  -13'd190,  13'd569,  13'd118,  -13'd861,  -13'd507,  13'd145,  -13'd377,  -13'd385,  13'd551,  -13'd164,  13'd328,  -13'd610,  
13'd292,  -13'd398,  13'd619,  13'd673,  -13'd802,  -13'd132,  -13'd167,  13'd805,  -13'd680,  -13'd648,  -13'd229,  13'd732,  13'd643,  13'd315,  13'd584,  13'd41,  
-13'd156,  13'd216,  -13'd827,  -13'd740,  -13'd374,  13'd694,  -13'd1254,  13'd172,  13'd728,  13'd66,  -13'd152,  13'd311,  -13'd318,  13'd47,  -13'd293,  13'd329,  
13'd169,  13'd662,  -13'd307,  13'd46,  13'd285,  13'd381,  13'd56,  -13'd12,  13'd217,  13'd438,  13'd284,  13'd892,  13'd300,  13'd185,  13'd106,  13'd388,  
13'd150,  -13'd442,  -13'd474,  13'd34,  -13'd375,  -13'd485,  13'd265,  13'd10,  13'd423,  -13'd303,  -13'd172,  -13'd399,  -13'd495,  13'd387,  -13'd201,  -13'd259,  
13'd577,  13'd341,  -13'd325,  13'd881,  13'd248,  -13'd1,  13'd132,  -13'd408,  -13'd141,  13'd463,  -13'd383,  -13'd383,  13'd635,  -13'd932,  13'd466,  -13'd115,  
13'd794,  -13'd72,  13'd296,  13'd37,  13'd134,  -13'd514,  -13'd722,  -13'd27,  
-13'd1040,  -13'd66,  -13'd714,  -13'd125,  -13'd307,  13'd335,  13'd314,  -13'd639,  13'd245,  13'd178,  13'd674,  -13'd388,  13'd388,  -13'd389,  13'd264,  -13'd402,  
-13'd461,  -13'd58,  -13'd18,  13'd853,  -13'd352,  -13'd317,  13'd392,  -13'd1006,  -13'd282,  13'd48,  13'd22,  13'd1027,  13'd363,  -13'd720,  13'd727,  -13'd40,  
13'd131,  -13'd310,  13'd143,  13'd40,  -13'd400,  -13'd3,  -13'd318,  13'd290,  13'd570,  13'd212,  -13'd607,  13'd791,  -13'd779,  13'd4,  13'd886,  -13'd320,  
13'd189,  13'd102,  13'd230,  13'd87,  -13'd59,  13'd109,  -13'd19,  -13'd357,  13'd743,  -13'd734,  13'd694,  -13'd874,  13'd383,  13'd628,  13'd232,  -13'd307,  
13'd66,  13'd264,  -13'd154,  -13'd65,  13'd187,  -13'd436,  13'd641,  13'd196,  -13'd6,  13'd440,  -13'd636,  13'd958,  -13'd538,  13'd870,  -13'd414,  13'd122,  
-13'd307,  13'd28,  13'd484,  13'd370,  -13'd40,  13'd556,  -13'd248,  13'd140,  -13'd45,  13'd426,  -13'd387,  13'd490,  -13'd579,  13'd395,  13'd399,  13'd118,  
-13'd356,  13'd680,  -13'd627,  13'd122,  13'd515,  -13'd266,  -13'd169,  -13'd232,  13'd645,  13'd12,  -13'd115,  13'd179,  -13'd191,  13'd762,  13'd358,  13'd206,  
-13'd7,  -13'd139,  -13'd281,  13'd886,  13'd120,  -13'd764,  13'd668,  -13'd764,  
-13'd307,  -13'd794,  13'd510,  13'd174,  -13'd778,  -13'd202,  -13'd11,  13'd908,  -13'd754,  -13'd556,  -13'd335,  -13'd250,  -13'd635,  -13'd51,  13'd39,  13'd331,  
-13'd171,  -13'd303,  -13'd467,  -13'd71,  -13'd371,  13'd202,  13'd351,  13'd119,  -13'd268,  13'd378,  13'd533,  13'd85,  -13'd542,  -13'd193,  -13'd652,  13'd405,  
13'd140,  13'd718,  -13'd166,  -13'd156,  13'd280,  -13'd92,  -13'd462,  -13'd195,  -13'd104,  13'd149,  13'd649,  -13'd543,  -13'd409,  -13'd469,  13'd308,  -13'd344,  
13'd448,  13'd331,  13'd209,  13'd42,  -13'd1065,  -13'd492,  13'd215,  -13'd503,  -13'd540,  13'd778,  13'd18,  -13'd391,  -13'd397,  13'd135,  13'd1386,  -13'd232,  
-13'd138,  -13'd987,  -13'd157,  -13'd555,  -13'd212,  -13'd25,  13'd737,  -13'd223,  -13'd264,  13'd161,  -13'd336,  -13'd58,  -13'd257,  13'd568,  13'd13,  13'd430,  
13'd25,  -13'd561,  13'd706,  13'd683,  -13'd332,  13'd448,  -13'd548,  -13'd643,  13'd657,  -13'd215,  -13'd114,  -13'd317,  -13'd306,  13'd65,  13'd414,  13'd217,  
13'd112,  13'd218,  -13'd36,  -13'd66,  13'd726,  13'd1011,  13'd244,  -13'd399,  13'd227,  13'd1103,  13'd440,  -13'd136,  -13'd241,  13'd1520,  -13'd603,  13'd108,  
13'd255,  -13'd859,  13'd543,  -13'd137,  -13'd616,  -13'd641,  -13'd285,  -13'd377,  
13'd242,  -13'd319,  13'd586,  13'd725,  -13'd229,  -13'd230,  -13'd355,  -13'd149,  -13'd83,  13'd828,  13'd224,  13'd114,  -13'd245,  13'd902,  13'd537,  13'd828,  
-13'd203,  13'd371,  13'd191,  -13'd670,  13'd701,  13'd255,  -13'd298,  13'd159,  -13'd706,  13'd121,  13'd186,  13'd270,  -13'd514,  13'd357,  13'd185,  13'd711,  
-13'd220,  13'd81,  13'd183,  -13'd207,  13'd192,  -13'd1164,  -13'd577,  13'd71,  -13'd913,  13'd460,  -13'd404,  -13'd405,  13'd895,  13'd435,  13'd297,  -13'd815,  
13'd280,  -13'd68,  -13'd51,  13'd67,  13'd225,  -13'd77,  -13'd491,  -13'd812,  -13'd394,  13'd483,  13'd230,  13'd891,  13'd428,  13'd89,  13'd368,  13'd546,  
13'd351,  13'd377,  13'd307,  -13'd797,  13'd424,  -13'd73,  13'd819,  13'd378,  -13'd249,  -13'd561,  -13'd651,  -13'd204,  13'd793,  -13'd358,  -13'd509,  13'd201,  
13'd589,  -13'd197,  13'd176,  13'd397,  13'd526,  13'd519,  -13'd423,  -13'd301,  -13'd110,  -13'd68,  -13'd213,  -13'd242,  -13'd582,  13'd216,  13'd271,  -13'd69,  
13'd549,  -13'd927,  -13'd292,  -13'd299,  -13'd48,  -13'd622,  13'd440,  -13'd1062,  -13'd46,  -13'd827,  -13'd270,  -13'd271,  13'd296,  -13'd74,  -13'd144,  13'd448,  
13'd179,  -13'd518,  -13'd416,  13'd395,  -13'd295,  -13'd809,  13'd320,  13'd94,  
13'd53,  13'd200,  -13'd483,  13'd470,  -13'd302,  13'd683,  13'd76,  -13'd412,  -13'd330,  -13'd755,  -13'd555,  -13'd516,  13'd272,  -13'd181,  -13'd557,  13'd401,  
-13'd156,  13'd183,  -13'd686,  13'd165,  -13'd455,  13'd82,  13'd503,  13'd158,  -13'd114,  13'd362,  -13'd505,  -13'd596,  -13'd173,  -13'd403,  -13'd512,  -13'd4,  
-13'd271,  13'd22,  13'd318,  -13'd467,  -13'd146,  13'd353,  -13'd441,  -13'd437,  13'd339,  -13'd25,  -13'd150,  13'd36,  -13'd305,  13'd129,  -13'd826,  -13'd26,  
13'd417,  -13'd732,  -13'd59,  -13'd540,  -13'd421,  -13'd122,  -13'd227,  -13'd37,  -13'd288,  13'd36,  -13'd605,  13'd67,  -13'd403,  -13'd153,  13'd798,  -13'd282,  
-13'd739,  -13'd657,  -13'd716,  -13'd143,  -13'd338,  -13'd179,  13'd509,  -13'd400,  -13'd377,  13'd155,  -13'd503,  13'd666,  -13'd282,  13'd75,  -13'd581,  13'd161,  
-13'd324,  13'd756,  -13'd110,  -13'd3,  -13'd329,  13'd91,  13'd223,  -13'd186,  13'd239,  -13'd629,  13'd507,  13'd574,  -13'd4,  13'd106,  13'd123,  13'd0,  
-13'd444,  -13'd655,  -13'd48,  -13'd603,  -13'd868,  -13'd34,  -13'd24,  13'd74,  -13'd797,  -13'd339,  -13'd674,  13'd256,  -13'd496,  -13'd146,  13'd99,  -13'd667,  
-13'd787,  13'd505,  -13'd520,  -13'd670,  -13'd59,  -13'd40,  13'd529,  13'd146,  
13'd471,  -13'd203,  -13'd705,  13'd275,  13'd310,  -13'd372,  13'd41,  13'd130,  -13'd284,  13'd281,  13'd602,  -13'd42,  13'd177,  -13'd375,  13'd195,  13'd18,  
-13'd768,  13'd188,  13'd110,  -13'd385,  -13'd137,  -13'd352,  -13'd517,  13'd235,  -13'd113,  -13'd231,  -13'd456,  13'd271,  -13'd201,  -13'd133,  -13'd199,  13'd183,  
13'd6,  -13'd509,  13'd9,  13'd437,  -13'd560,  -13'd148,  13'd92,  -13'd99,  -13'd123,  -13'd263,  -13'd435,  -13'd369,  13'd102,  -13'd183,  -13'd581,  -13'd403,  
-13'd132,  -13'd122,  -13'd408,  -13'd25,  -13'd178,  -13'd294,  13'd355,  13'd117,  13'd54,  -13'd181,  -13'd322,  13'd510,  13'd38,  -13'd431,  13'd425,  -13'd156,  
13'd459,  -13'd939,  13'd64,  -13'd259,  13'd244,  -13'd328,  13'd183,  -13'd357,  -13'd144,  13'd466,  -13'd462,  13'd303,  -13'd37,  -13'd17,  -13'd275,  13'd343,  
-13'd147,  13'd396,  13'd402,  -13'd764,  -13'd616,  -13'd113,  -13'd459,  13'd409,  -13'd11,  -13'd742,  13'd378,  -13'd294,  13'd288,  -13'd58,  13'd594,  -13'd298,  
-13'd432,  -13'd476,  13'd53,  13'd357,  13'd139,  13'd115,  -13'd885,  -13'd526,  -13'd38,  -13'd581,  -13'd257,  -13'd697,  -13'd395,  -13'd169,  13'd117,  -13'd407,  
13'd82,  13'd25,  -13'd659,  -13'd639,  -13'd622,  -13'd394,  -13'd415,  -13'd8,  
-13'd140,  13'd150,  -13'd432,  13'd1,  -13'd518,  13'd588,  13'd143,  13'd80,  -13'd75,  -13'd817,  13'd537,  -13'd126,  -13'd321,  13'd433,  -13'd432,  -13'd82,  
-13'd319,  -13'd403,  -13'd898,  -13'd508,  -13'd403,  -13'd727,  -13'd86,  -13'd118,  -13'd151,  -13'd590,  -13'd493,  -13'd685,  -13'd230,  13'd388,  -13'd176,  -13'd552,  
-13'd197,  -13'd572,  13'd84,  -13'd56,  13'd702,  -13'd562,  -13'd50,  -13'd636,  -13'd693,  -13'd833,  -13'd132,  -13'd296,  -13'd498,  13'd108,  -13'd342,  -13'd125,  
13'd454,  13'd100,  -13'd410,  -13'd645,  13'd104,  13'd194,  -13'd935,  13'd489,  13'd225,  13'd230,  -13'd277,  -13'd222,  -13'd55,  -13'd144,  -13'd63,  -13'd102,  
13'd543,  -13'd561,  -13'd111,  -13'd681,  -13'd338,  -13'd62,  13'd378,  -13'd177,  -13'd218,  -13'd363,  -13'd416,  -13'd393,  -13'd295,  -13'd660,  -13'd406,  -13'd555,  
-13'd509,  -13'd570,  13'd22,  -13'd291,  13'd300,  -13'd392,  13'd80,  13'd90,  -13'd135,  13'd8,  -13'd148,  13'd153,  13'd155,  -13'd165,  13'd52,  -13'd82,  
-13'd1005,  -13'd576,  13'd577,  -13'd851,  -13'd442,  -13'd228,  -13'd371,  13'd536,  13'd121,  13'd122,  -13'd73,  -13'd439,  13'd136,  -13'd573,  -13'd527,  -13'd348,  
13'd133,  13'd112,  13'd98,  13'd57,  -13'd103,  13'd198,  13'd142,  -13'd137,  
13'd221,  -13'd283,  -13'd623,  13'd183,  13'd55,  13'd781,  -13'd42,  -13'd133,  -13'd55,  -13'd543,  -13'd1,  13'd57,  -13'd660,  -13'd664,  13'd603,  -13'd312,  
13'd181,  13'd501,  13'd161,  -13'd199,  13'd473,  13'd270,  -13'd469,  -13'd150,  -13'd256,  13'd290,  13'd413,  -13'd297,  -13'd302,  -13'd247,  -13'd284,  13'd231,  
-13'd69,  13'd88,  -13'd420,  -13'd609,  13'd217,  -13'd62,  13'd469,  -13'd175,  -13'd62,  -13'd682,  -13'd264,  -13'd387,  -13'd225,  -13'd80,  -13'd552,  -13'd181,  
13'd373,  13'd41,  -13'd491,  13'd600,  13'd615,  13'd205,  13'd763,  -13'd329,  13'd97,  13'd72,  -13'd359,  -13'd51,  13'd259,  -13'd56,  13'd228,  13'd13,  
-13'd490,  -13'd756,  13'd154,  -13'd730,  -13'd82,  -13'd348,  -13'd140,  -13'd622,  13'd476,  -13'd181,  13'd566,  -13'd426,  13'd455,  13'd476,  -13'd215,  -13'd41,  
13'd247,  13'd592,  13'd30,  -13'd7,  13'd77,  -13'd787,  13'd153,  -13'd338,  13'd197,  13'd292,  -13'd826,  -13'd318,  -13'd90,  -13'd26,  -13'd424,  -13'd217,  
-13'd196,  -13'd343,  -13'd630,  13'd247,  -13'd132,  -13'd291,  -13'd756,  -13'd156,  -13'd665,  13'd359,  -13'd285,  -13'd271,  -13'd317,  -13'd88,  -13'd534,  -13'd395,  
-13'd306,  -13'd355,  13'd422,  -13'd281,  13'd104,  -13'd82,  -13'd137,  -13'd585,  
-13'd377,  -13'd315,  13'd233,  13'd251,  -13'd977,  13'd544,  13'd276,  -13'd33,  13'd372,  -13'd111,  -13'd444,  13'd372,  -13'd19,  13'd576,  13'd744,  -13'd221,  
-13'd1370,  -13'd295,  13'd807,  -13'd563,  13'd39,  -13'd649,  13'd411,  13'd17,  13'd302,  -13'd139,  13'd1108,  -13'd421,  -13'd1262,  13'd275,  -13'd120,  -13'd146,  
-13'd403,  13'd570,  -13'd1176,  -13'd366,  13'd165,  13'd1003,  13'd875,  -13'd106,  13'd409,  -13'd321,  -13'd336,  -13'd407,  -13'd13,  13'd45,  -13'd104,  13'd367,  
-13'd441,  13'd416,  13'd475,  13'd96,  13'd99,  13'd45,  13'd150,  -13'd179,  13'd496,  13'd606,  13'd44,  -13'd125,  -13'd1209,  -13'd0,  13'd889,  -13'd282,  
13'd124,  -13'd747,  13'd493,  13'd281,  13'd694,  -13'd545,  13'd1702,  -13'd39,  -13'd858,  13'd137,  -13'd38,  13'd78,  -13'd134,  -13'd390,  -13'd878,  -13'd674,  
13'd286,  13'd334,  13'd117,  -13'd14,  13'd493,  -13'd557,  -13'd409,  -13'd321,  13'd112,  13'd951,  13'd264,  13'd88,  13'd74,  13'd231,  -13'd685,  13'd258,  
13'd495,  -13'd363,  13'd1061,  13'd756,  13'd431,  -13'd303,  -13'd692,  13'd669,  13'd413,  13'd955,  -13'd531,  -13'd1012,  -13'd367,  13'd47,  -13'd60,  -13'd147,  
13'd454,  13'd313,  13'd785,  13'd715,  -13'd642,  13'd540,  13'd694,  13'd479,  
-13'd669,  -13'd553,  13'd468,  13'd187,  -13'd493,  -13'd832,  -13'd472,  -13'd209,  13'd233,  13'd192,  -13'd227,  13'd426,  13'd30,  -13'd766,  13'd303,  13'd19,  
-13'd174,  -13'd431,  -13'd684,  -13'd608,  -13'd445,  -13'd132,  -13'd233,  -13'd412,  13'd250,  -13'd41,  -13'd300,  13'd67,  -13'd125,  13'd164,  13'd689,  13'd510,  
13'd226,  -13'd300,  -13'd366,  13'd161,  -13'd68,  13'd219,  13'd54,  -13'd150,  -13'd73,  13'd199,  -13'd914,  13'd287,  13'd171,  13'd351,  -13'd107,  -13'd62,  
-13'd300,  13'd386,  -13'd71,  -13'd361,  -13'd308,  13'd354,  -13'd75,  -13'd427,  -13'd573,  13'd50,  -13'd283,  -13'd471,  -13'd118,  -13'd225,  -13'd105,  13'd409,  
-13'd12,  -13'd699,  13'd253,  -13'd81,  -13'd446,  13'd138,  -13'd343,  -13'd51,  13'd313,  -13'd463,  -13'd106,  -13'd198,  13'd115,  13'd24,  -13'd48,  13'd78,  
-13'd74,  -13'd249,  -13'd219,  -13'd511,  -13'd54,  13'd340,  13'd26,  -13'd855,  13'd426,  13'd72,  -13'd81,  13'd281,  -13'd420,  -13'd517,  13'd132,  -13'd160,  
13'd361,  13'd62,  -13'd337,  -13'd195,  -13'd588,  -13'd73,  -13'd349,  13'd145,  -13'd43,  -13'd18,  -13'd365,  -13'd901,  -13'd212,  13'd170,  13'd73,  13'd45,  
-13'd36,  13'd181,  -13'd263,  -13'd128,  -13'd279,  13'd580,  -13'd264,  13'd187,  
13'd1174,  13'd86,  13'd226,  -13'd27,  -13'd245,  13'd196,  13'd204,  -13'd678,  13'd587,  -13'd2,  13'd246,  -13'd883,  13'd12,  -13'd590,  -13'd328,  13'd414,  
13'd321,  -13'd280,  13'd154,  13'd208,  13'd346,  13'd610,  13'd87,  13'd924,  13'd324,  13'd468,  13'd15,  13'd417,  -13'd361,  13'd602,  13'd363,  13'd255,  
13'd247,  -13'd508,  13'd423,  13'd558,  13'd21,  13'd656,  13'd794,  -13'd807,  -13'd296,  13'd731,  -13'd729,  -13'd442,  13'd159,  -13'd633,  -13'd789,  -13'd702,  
-13'd157,  -13'd178,  13'd439,  -13'd597,  13'd235,  13'd258,  13'd277,  -13'd123,  -13'd623,  13'd339,  13'd395,  13'd206,  -13'd405,  -13'd61,  -13'd510,  13'd7,  
13'd702,  -13'd1044,  13'd688,  13'd229,  -13'd69,  13'd884,  -13'd279,  -13'd475,  -13'd456,  -13'd698,  13'd27,  -13'd866,  -13'd141,  -13'd292,  13'd737,  -13'd190,  
-13'd205,  13'd169,  13'd588,  -13'd15,  -13'd894,  -13'd607,  13'd300,  -13'd454,  -13'd214,  13'd458,  13'd495,  13'd369,  13'd744,  13'd340,  13'd512,  13'd605,  
13'd510,  13'd907,  -13'd696,  -13'd24,  -13'd80,  -13'd541,  13'd381,  13'd1443,  13'd73,  -13'd527,  13'd72,  -13'd532,  13'd45,  13'd991,  -13'd552,  13'd169,  
13'd115,  -13'd735,  -13'd492,  -13'd695,  13'd515,  -13'd442,  -13'd329,  -13'd119,  
-13'd732,  -13'd328,  -13'd508,  13'd109,  13'd36,  13'd252,  13'd2,  -13'd28,  -13'd375,  -13'd215,  13'd347,  13'd53,  -13'd406,  13'd473,  -13'd235,  13'd115,  
-13'd431,  -13'd209,  -13'd343,  -13'd6,  13'd551,  -13'd36,  -13'd184,  -13'd129,  13'd128,  13'd120,  13'd488,  13'd491,  13'd320,  -13'd428,  -13'd120,  -13'd1137,  
-13'd135,  13'd54,  13'd451,  -13'd337,  13'd312,  13'd188,  -13'd665,  13'd158,  -13'd260,  13'd615,  -13'd80,  13'd33,  -13'd954,  13'd485,  -13'd261,  13'd180,  
13'd427,  -13'd197,  13'd112,  13'd114,  -13'd431,  13'd771,  13'd932,  -13'd106,  13'd233,  -13'd222,  13'd649,  -13'd718,  13'd70,  13'd722,  13'd858,  -13'd501,  
-13'd524,  -13'd30,  13'd135,  -13'd23,  13'd348,  -13'd440,  -13'd207,  -13'd50,  13'd384,  -13'd300,  -13'd617,  13'd139,  -13'd728,  -13'd226,  -13'd557,  13'd262,  
-13'd277,  13'd164,  13'd16,  -13'd530,  13'd177,  13'd434,  13'd173,  -13'd37,  -13'd8,  13'd455,  13'd217,  13'd806,  -13'd827,  -13'd239,  13'd77,  13'd534,  
-13'd235,  13'd284,  -13'd112,  13'd319,  13'd187,  13'd93,  -13'd484,  13'd49,  13'd71,  -13'd26,  -13'd29,  13'd86,  -13'd34,  13'd33,  13'd205,  -13'd940,  
13'd498,  -13'd96,  13'd552,  -13'd229,  13'd700,  13'd434,  13'd224,  13'd195,  
13'd183,  13'd132,  -13'd571,  -13'd86,  13'd1180,  -13'd19,  13'd244,  13'd1090,  -13'd65,  -13'd208,  13'd370,  13'd594,  -13'd375,  -13'd705,  -13'd237,  -13'd486,  
13'd1048,  13'd512,  -13'd483,  13'd216,  13'd180,  -13'd25,  -13'd83,  13'd91,  13'd40,  13'd707,  -13'd311,  13'd6,  -13'd470,  13'd548,  13'd324,  -13'd637,  
13'd213,  -13'd255,  -13'd314,  13'd115,  -13'd2,  -13'd228,  13'd138,  13'd333,  -13'd257,  -13'd365,  13'd916,  -13'd272,  -13'd152,  13'd634,  -13'd399,  13'd279,  
-13'd115,  13'd652,  13'd210,  13'd669,  13'd330,  13'd40,  -13'd375,  -13'd170,  -13'd447,  -13'd200,  -13'd319,  13'd440,  -13'd80,  13'd83,  -13'd121,  13'd320,  
13'd383,  13'd558,  -13'd353,  13'd329,  13'd430,  13'd508,  -13'd380,  13'd173,  13'd356,  13'd189,  13'd388,  -13'd224,  -13'd153,  13'd400,  -13'd464,  13'd227,  
-13'd666,  13'd323,  -13'd363,  13'd1110,  13'd526,  -13'd525,  -13'd500,  -13'd432,  -13'd228,  13'd560,  -13'd827,  -13'd232,  13'd334,  13'd675,  -13'd70,  -13'd391,  
13'd220,  -13'd332,  -13'd467,  13'd598,  13'd91,  -13'd569,  -13'd427,  13'd534,  13'd461,  -13'd379,  -13'd631,  13'd674,  -13'd139,  -13'd1067,  -13'd10,  -13'd424,  
-13'd252,  13'd990,  -13'd512,  13'd526,  -13'd211,  13'd98,  -13'd99,  -13'd338,  
13'd677,  13'd8,  -13'd349,  13'd171,  -13'd97,  13'd358,  -13'd517,  13'd747,  -13'd276,  -13'd137,  -13'd184,  -13'd591,  -13'd344,  -13'd369,  -13'd648,  13'd708,  
13'd180,  -13'd612,  -13'd145,  -13'd244,  13'd657,  13'd247,  -13'd423,  -13'd299,  -13'd466,  13'd314,  -13'd579,  -13'd238,  -13'd760,  -13'd413,  13'd346,  -13'd358,  
-13'd24,  13'd103,  -13'd0,  -13'd0,  13'd275,  13'd256,  -13'd259,  13'd134,  13'd115,  13'd58,  -13'd521,  13'd150,  -13'd220,  13'd347,  -13'd88,  13'd32,  
-13'd426,  -13'd165,  13'd66,  -13'd239,  -13'd535,  -13'd411,  -13'd579,  -13'd366,  -13'd250,  13'd14,  13'd344,  -13'd330,  13'd301,  13'd608,  -13'd250,  -13'd26,  
-13'd266,  13'd489,  13'd170,  13'd409,  -13'd445,  -13'd54,  13'd424,  -13'd146,  13'd32,  13'd374,  -13'd133,  13'd515,  -13'd106,  13'd212,  -13'd417,  13'd350,  
-13'd625,  -13'd96,  -13'd135,  13'd239,  13'd253,  -13'd371,  -13'd578,  13'd238,  -13'd114,  -13'd298,  -13'd303,  -13'd313,  -13'd18,  -13'd518,  13'd469,  -13'd170,  
13'd278,  13'd35,  -13'd202,  -13'd174,  -13'd0,  -13'd185,  13'd438,  13'd680,  -13'd39,  -13'd715,  -13'd323,  13'd209,  13'd381,  13'd214,  -13'd223,  -13'd216,  
13'd98,  13'd571,  13'd568,  13'd47,  13'd162,  13'd390,  -13'd109,  13'd704,  
13'd1172,  13'd88,  -13'd23,  13'd555,  13'd665,  13'd21,  -13'd117,  13'd340,  -13'd726,  -13'd282,  -13'd53,  -13'd544,  13'd6,  -13'd106,  13'd330,  13'd241,  
13'd254,  13'd413,  -13'd786,  13'd448,  -13'd664,  13'd37,  13'd260,  13'd879,  -13'd580,  13'd748,  13'd234,  13'd680,  -13'd581,  13'd293,  -13'd46,  -13'd413,  
-13'd86,  -13'd354,  13'd104,  -13'd141,  13'd423,  13'd507,  13'd871,  -13'd24,  13'd682,  -13'd103,  -13'd605,  -13'd817,  -13'd526,  -13'd101,  -13'd685,  13'd245,  
-13'd126,  13'd71,  -13'd584,  -13'd472,  13'd692,  13'd230,  -13'd192,  -13'd499,  13'd807,  13'd879,  -13'd71,  -13'd176,  13'd397,  13'd12,  -13'd850,  13'd2,  
13'd59,  13'd678,  13'd669,  13'd374,  13'd500,  13'd268,  13'd35,  -13'd122,  -13'd243,  13'd962,  -13'd355,  -13'd272,  13'd770,  13'd625,  -13'd96,  13'd162,  
-13'd605,  13'd549,  -13'd153,  13'd53,  -13'd240,  13'd381,  -13'd280,  -13'd15,  -13'd19,  13'd691,  -13'd97,  13'd517,  13'd907,  -13'd176,  13'd314,  -13'd220,  
13'd105,  -13'd71,  -13'd246,  13'd303,  -13'd548,  13'd178,  13'd723,  13'd692,  -13'd774,  -13'd17,  13'd165,  13'd171,  13'd258,  -13'd234,  13'd744,  13'd445,  
-13'd625,  13'd272,  13'd187,  -13'd161,  -13'd239,  13'd92,  13'd81,  13'd915,  
-13'd1121,  -13'd378,  13'd566,  13'd36,  -13'd315,  -13'd527,  13'd293,  13'd1088,  13'd110,  13'd122,  -13'd358,  13'd1119,  -13'd15,  13'd408,  13'd877,  -13'd515,  
-13'd154,  13'd538,  13'd198,  -13'd685,  13'd205,  -13'd836,  13'd9,  -13'd160,  -13'd233,  -13'd494,  13'd863,  -13'd96,  -13'd14,  13'd735,  -13'd179,  -13'd137,  
-13'd576,  -13'd283,  -13'd193,  13'd175,  -13'd204,  -13'd584,  13'd87,  13'd351,  13'd52,  -13'd478,  13'd726,  13'd225,  13'd209,  13'd155,  13'd100,  13'd1009,  
-13'd729,  13'd500,  13'd974,  -13'd1373,  -13'd403,  -13'd1104,  -13'd610,  13'd358,  -13'd384,  -13'd242,  13'd473,  13'd73,  -13'd402,  13'd15,  13'd39,  13'd292,  
-13'd1232,  13'd467,  13'd327,  -13'd712,  13'd196,  -13'd1266,  -13'd141,  13'd156,  -13'd48,  -13'd586,  -13'd37,  -13'd229,  13'd1126,  -13'd127,  -13'd506,  -13'd98,  
13'd52,  13'd661,  -13'd151,  -13'd533,  -13'd109,  13'd357,  13'd90,  13'd199,  -13'd238,  13'd349,  -13'd334,  13'd641,  13'd116,  -13'd64,  13'd106,  13'd181,  
13'd455,  13'd24,  -13'd111,  -13'd237,  -13'd158,  -13'd1204,  -13'd84,  -13'd414,  13'd64,  -13'd735,  -13'd796,  -13'd16,  13'd389,  13'd100,  13'd497,  -13'd198,  
13'd403,  13'd354,  -13'd54,  13'd273,  -13'd21,  13'd87,  -13'd706,  13'd935,  
13'd280,  13'd5,  13'd716,  -13'd314,  -13'd416,  13'd83,  13'd580,  -13'd463,  13'd951,  13'd392,  13'd166,  13'd225,  -13'd56,  -13'd771,  -13'd479,  13'd867,  
13'd441,  13'd7,  13'd732,  13'd413,  -13'd214,  13'd513,  13'd114,  13'd521,  13'd426,  13'd396,  -13'd37,  -13'd234,  -13'd609,  -13'd228,  -13'd969,  -13'd958,  
13'd608,  -13'd310,  -13'd113,  -13'd86,  -13'd591,  13'd838,  13'd954,  -13'd584,  13'd446,  -13'd43,  13'd111,  13'd330,  -13'd535,  -13'd48,  13'd58,  -13'd249,  
13'd201,  -13'd772,  13'd32,  -13'd620,  13'd129,  -13'd131,  13'd67,  13'd210,  -13'd928,  13'd51,  13'd84,  -13'd307,  -13'd294,  -13'd242,  -13'd789,  -13'd285,  
13'd1217,  -13'd721,  -13'd211,  13'd460,  13'd931,  13'd409,  -13'd635,  13'd636,  -13'd28,  -13'd117,  13'd528,  13'd493,  -13'd747,  -13'd263,  13'd90,  13'd392,  
-13'd511,  13'd3,  -13'd376,  13'd140,  -13'd343,  13'd211,  -13'd350,  13'd915,  13'd285,  13'd331,  -13'd365,  13'd217,  13'd394,  13'd134,  13'd269,  -13'd250,  
-13'd208,  -13'd265,  -13'd378,  -13'd34,  -13'd663,  -13'd102,  13'd148,  13'd679,  -13'd300,  13'd225,  13'd104,  -13'd717,  13'd547,  13'd177,  13'd250,  -13'd215,  
-13'd607,  -13'd267,  -13'd469,  13'd45,  13'd378,  13'd266,  13'd22,  13'd459,  
13'd269,  -13'd27,  -13'd892,  13'd174,  -13'd695,  13'd197,  13'd136,  13'd343,  -13'd704,  -13'd213,  -13'd196,  13'd40,  -13'd273,  13'd254,  13'd229,  13'd893,  
13'd352,  -13'd338,  13'd512,  -13'd420,  -13'd478,  -13'd475,  -13'd236,  -13'd478,  13'd247,  -13'd750,  13'd137,  13'd150,  -13'd19,  13'd299,  -13'd122,  -13'd753,  
-13'd676,  13'd18,  -13'd693,  13'd293,  13'd478,  -13'd367,  -13'd531,  13'd236,  -13'd674,  -13'd909,  13'd19,  -13'd80,  13'd405,  -13'd70,  -13'd94,  13'd506,  
13'd483,  -13'd1111,  13'd195,  -13'd445,  -13'd347,  -13'd536,  13'd159,  13'd271,  -13'd532,  13'd203,  -13'd21,  13'd282,  -13'd28,  -13'd830,  -13'd816,  -13'd60,  
13'd547,  -13'd237,  13'd352,  13'd30,  -13'd566,  13'd86,  13'd398,  -13'd156,  13'd16,  13'd866,  -13'd709,  -13'd604,  13'd358,  -13'd236,  -13'd741,  -13'd26,  
-13'd165,  -13'd495,  13'd558,  -13'd534,  -13'd654,  13'd373,  13'd23,  13'd613,  -13'd836,  -13'd116,  -13'd390,  -13'd300,  13'd454,  -13'd124,  -13'd94,  13'd584,  
13'd226,  -13'd670,  13'd655,  -13'd585,  -13'd124,  -13'd1236,  -13'd458,  13'd139,  -13'd125,  -13'd398,  -13'd405,  -13'd261,  13'd163,  13'd374,  -13'd538,  13'd783,  
13'd572,  -13'd225,  13'd391,  -13'd345,  13'd247,  13'd5,  13'd599,  13'd915,  
-13'd474,  -13'd190,  -13'd534,  13'd70,  -13'd390,  -13'd541,  13'd158,  13'd22,  13'd320,  -13'd538,  -13'd389,  13'd314,  13'd81,  -13'd80,  13'd451,  -13'd359,  
-13'd147,  -13'd66,  13'd53,  13'd303,  13'd546,  13'd203,  -13'd24,  13'd37,  -13'd107,  -13'd321,  -13'd35,  -13'd596,  13'd239,  -13'd760,  -13'd354,  -13'd270,  
13'd559,  -13'd867,  -13'd888,  13'd450,  -13'd309,  -13'd805,  -13'd51,  -13'd622,  -13'd134,  13'd453,  -13'd334,  -13'd527,  -13'd452,  13'd20,  -13'd533,  13'd13,  
13'd324,  13'd310,  -13'd366,  -13'd156,  -13'd196,  13'd135,  13'd72,  -13'd251,  13'd405,  13'd132,  13'd110,  -13'd317,  -13'd587,  13'd30,  -13'd125,  13'd574,  
13'd143,  13'd6,  -13'd301,  -13'd93,  -13'd88,  -13'd3,  -13'd58,  13'd116,  13'd23,  -13'd240,  -13'd467,  13'd290,  -13'd336,  -13'd460,  -13'd374,  13'd434,  
13'd493,  -13'd452,  -13'd422,  13'd791,  -13'd511,  13'd287,  -13'd466,  -13'd405,  13'd418,  -13'd613,  13'd166,  -13'd824,  -13'd324,  -13'd4,  -13'd720,  13'd36,  
13'd378,  -13'd486,  -13'd247,  13'd32,  -13'd259,  13'd433,  13'd279,  13'd212,  13'd392,  -13'd147,  13'd342,  13'd118,  13'd424,  -13'd782,  -13'd67,  13'd107,  
-13'd289,  -13'd365,  -13'd195,  -13'd155,  -13'd505,  -13'd182,  13'd453,  -13'd10,  
13'd100,  -13'd389,  -13'd584,  13'd5,  -13'd116,  13'd166,  -13'd178,  -13'd598,  13'd520,  -13'd428,  13'd495,  -13'd408,  13'd327,  -13'd699,  -13'd174,  13'd127,  
-13'd177,  13'd309,  -13'd50,  13'd108,  13'd265,  13'd386,  13'd475,  13'd163,  13'd743,  13'd276,  13'd178,  -13'd189,  -13'd781,  -13'd178,  13'd475,  13'd351,  
13'd890,  13'd441,  13'd112,  -13'd136,  -13'd30,  13'd110,  13'd473,  -13'd407,  13'd464,  13'd596,  -13'd274,  13'd751,  -13'd151,  -13'd586,  -13'd753,  -13'd965,  
-13'd91,  -13'd374,  -13'd222,  13'd908,  13'd258,  13'd139,  13'd695,  13'd359,  -13'd541,  13'd725,  13'd216,  13'd39,  13'd357,  13'd504,  13'd67,  13'd34,  
13'd157,  -13'd710,  13'd183,  13'd1472,  13'd186,  13'd85,  13'd214,  13'd547,  13'd758,  -13'd560,  13'd124,  13'd133,  -13'd901,  13'd278,  -13'd477,  -13'd514,  
13'd746,  13'd495,  -13'd243,  -13'd14,  13'd611,  13'd37,  13'd778,  -13'd22,  13'd279,  -13'd419,  13'd249,  -13'd176,  13'd441,  -13'd34,  -13'd276,  13'd550,  
13'd493,  13'd611,  -13'd545,  -13'd166,  -13'd426,  13'd204,  -13'd143,  13'd716,  -13'd795,  13'd73,  13'd299,  -13'd1303,  13'd46,  13'd833,  13'd42,  13'd267,  
-13'd278,  -13'd276,  -13'd221,  -13'd151,  13'd458,  -13'd132,  13'd559,  13'd325,  
13'd418,  -13'd205,  13'd368,  -13'd221,  -13'd703,  -13'd206,  13'd284,  13'd405,  13'd71,  -13'd60,  -13'd234,  -13'd257,  -13'd155,  -13'd293,  13'd167,  13'd709,  
-13'd503,  -13'd565,  -13'd323,  -13'd478,  13'd43,  13'd285,  -13'd237,  -13'd141,  13'd8,  13'd97,  -13'd719,  -13'd187,  13'd824,  -13'd478,  -13'd69,  13'd803,  
-13'd244,  13'd530,  -13'd32,  13'd185,  -13'd217,  -13'd420,  -13'd752,  13'd71,  13'd37,  13'd275,  13'd907,  13'd178,  13'd0,  -13'd320,  13'd398,  -13'd306,  
13'd534,  13'd807,  13'd357,  -13'd37,  -13'd338,  -13'd722,  13'd1059,  -13'd745,  -13'd4,  13'd628,  13'd380,  -13'd753,  -13'd550,  13'd202,  -13'd263,  -13'd2,  
13'd496,  13'd449,  13'd110,  13'd236,  -13'd10,  -13'd1115,  -13'd539,  13'd421,  13'd584,  -13'd1117,  13'd737,  -13'd943,  -13'd969,  -13'd463,  -13'd78,  13'd96,  
-13'd59,  13'd470,  13'd180,  -13'd315,  13'd444,  13'd638,  -13'd465,  -13'd162,  13'd232,  13'd121,  -13'd419,  13'd53,  13'd331,  13'd467,  -13'd790,  13'd77,  
13'd239,  13'd907,  -13'd345,  -13'd1114,  13'd951,  -13'd526,  -13'd881,  -13'd405,  13'd537,  -13'd371,  13'd133,  -13'd171,  13'd259,  13'd107,  13'd490,  -13'd9,  
-13'd376,  13'd478,  13'd619,  13'd446,  13'd525,  13'd739,  13'd276,  -13'd485,  
-13'd895,  13'd255,  -13'd202,  13'd197,  13'd24,  -13'd261,  13'd567,  -13'd816,  -13'd949,  13'd0,  13'd352,  13'd826,  13'd45,  13'd59,  -13'd22,  13'd232,  
-13'd713,  13'd102,  13'd431,  -13'd81,  -13'd246,  -13'd188,  13'd417,  13'd15,  13'd395,  -13'd917,  -13'd18,  13'd127,  13'd554,  -13'd191,  13'd576,  -13'd113,  
13'd160,  -13'd380,  13'd460,  13'd122,  -13'd834,  13'd83,  13'd480,  13'd653,  -13'd162,  -13'd348,  -13'd379,  -13'd695,  13'd200,  13'd173,  13'd454,  -13'd158,  
-13'd133,  -13'd726,  -13'd487,  13'd396,  -13'd347,  13'd99,  13'd434,  13'd237,  13'd326,  13'd46,  13'd560,  13'd275,  -13'd70,  13'd489,  -13'd64,  -13'd392,  
13'd656,  13'd789,  13'd370,  13'd782,  13'd126,  -13'd700,  -13'd35,  13'd98,  13'd32,  -13'd396,  13'd171,  13'd679,  13'd304,  13'd27,  13'd470,  13'd628,  
13'd324,  13'd227,  13'd241,  -13'd618,  -13'd555,  13'd634,  13'd510,  13'd173,  -13'd279,  13'd594,  13'd60,  13'd131,  -13'd828,  -13'd450,  13'd145,  -13'd34,  
13'd63,  -13'd204,  13'd896,  -13'd540,  13'd165,  13'd274,  -13'd278,  -13'd621,  -13'd111,  13'd590,  13'd172,  -13'd389,  -13'd219,  13'd1034,  -13'd359,  -13'd449,  
13'd34,  -13'd926,  13'd349,  13'd150,  13'd430,  13'd473,  13'd874,  13'd607,  
13'd172,  13'd107,  13'd358,  13'd115,  -13'd146,  13'd83,  13'd559,  13'd173,  13'd107,  13'd98,  -13'd335,  13'd169,  13'd447,  13'd178,  -13'd376,  -13'd221,  
-13'd67,  -13'd957,  -13'd78,  -13'd394,  -13'd706,  13'd119,  13'd126,  13'd7,  -13'd153,  -13'd600,  13'd82,  -13'd755,  -13'd539,  13'd229,  13'd564,  -13'd116,  
13'd68,  -13'd630,  -13'd509,  -13'd185,  13'd695,  -13'd546,  -13'd620,  -13'd12,  -13'd411,  13'd48,  13'd381,  -13'd411,  13'd497,  13'd126,  -13'd771,  -13'd644,  
13'd11,  -13'd879,  -13'd802,  13'd242,  13'd200,  -13'd315,  -13'd472,  13'd592,  13'd67,  13'd0,  13'd70,  -13'd343,  -13'd420,  13'd23,  -13'd263,  -13'd604,  
-13'd349,  -13'd97,  -13'd247,  13'd489,  -13'd992,  -13'd199,  -13'd99,  -13'd481,  -13'd485,  -13'd21,  -13'd459,  13'd284,  13'd304,  13'd281,  13'd444,  13'd292,  
-13'd397,  13'd411,  -13'd458,  13'd247,  -13'd852,  -13'd246,  -13'd492,  13'd247,  13'd183,  -13'd221,  -13'd382,  13'd149,  -13'd318,  -13'd220,  -13'd263,  -13'd907,  
-13'd58,  -13'd411,  -13'd114,  -13'd398,  -13'd416,  13'd140,  -13'd749,  -13'd507,  13'd348,  -13'd292,  -13'd403,  13'd424,  13'd257,  13'd555,  -13'd192,  13'd164,  
-13'd25,  13'd174,  13'd197,  13'd23,  13'd582,  13'd308,  -13'd401,  13'd80,  
-13'd661,  -13'd481,  -13'd16,  13'd159,  -13'd350,  -13'd271,  -13'd58,  -13'd213,  13'd510,  -13'd408,  13'd591,  13'd52,  -13'd183,  -13'd277,  13'd514,  -13'd312,  
13'd146,  -13'd164,  -13'd516,  -13'd864,  -13'd250,  -13'd760,  -13'd508,  -13'd899,  -13'd420,  -13'd364,  -13'd89,  -13'd334,  -13'd284,  -13'd704,  -13'd89,  -13'd522,  
-13'd76,  -13'd263,  -13'd26,  -13'd152,  -13'd427,  13'd32,  -13'd74,  -13'd172,  13'd380,  13'd333,  -13'd214,  13'd130,  -13'd460,  -13'd311,  -13'd536,  -13'd112,  
-13'd300,  -13'd777,  13'd22,  13'd12,  -13'd495,  -13'd400,  13'd467,  13'd671,  -13'd85,  13'd648,  13'd207,  -13'd777,  -13'd529,  -13'd469,  -13'd617,  -13'd287,  
-13'd394,  -13'd574,  13'd36,  13'd140,  13'd352,  13'd491,  -13'd67,  -13'd446,  -13'd669,  13'd416,  13'd25,  13'd486,  13'd313,  13'd337,  -13'd513,  -13'd950,  
13'd243,  13'd363,  -13'd658,  13'd307,  -13'd104,  13'd70,  -13'd49,  -13'd819,  -13'd432,  13'd277,  13'd201,  -13'd165,  13'd174,  -13'd830,  13'd317,  13'd283,  
13'd649,  -13'd469,  13'd308,  -13'd408,  -13'd73,  -13'd742,  -13'd367,  -13'd258,  -13'd554,  13'd639,  -13'd93,  -13'd690,  -13'd527,  13'd536,  13'd72,  13'd247,  
-13'd278,  -13'd959,  13'd375,  13'd372,  -13'd688,  -13'd604,  -13'd103,  -13'd295,  
-13'd725,  -13'd95,  -13'd741,  -13'd304,  -13'd675,  -13'd123,  -13'd504,  13'd180,  13'd487,  -13'd527,  13'd193,  13'd69,  -13'd499,  -13'd19,  13'd43,  -13'd870,  
-13'd100,  13'd364,  -13'd871,  13'd190,  -13'd473,  13'd391,  13'd155,  -13'd22,  -13'd177,  13'd446,  13'd350,  13'd48,  13'd91,  13'd406,  13'd826,  -13'd398,  
13'd769,  -13'd77,  -13'd324,  -13'd351,  -13'd123,  -13'd223,  -13'd290,  13'd136,  13'd531,  13'd104,  13'd872,  13'd287,  13'd548,  13'd294,  13'd477,  13'd219,  
-13'd102,  13'd169,  13'd806,  13'd565,  -13'd845,  -13'd69,  13'd32,  -13'd684,  13'd235,  13'd104,  -13'd168,  -13'd148,  -13'd630,  13'd501,  13'd305,  13'd132,  
-13'd587,  13'd202,  -13'd382,  -13'd256,  13'd192,  -13'd480,  13'd21,  -13'd374,  13'd345,  -13'd1113,  -13'd137,  -13'd244,  -13'd992,  13'd1014,  -13'd368,  13'd798,  
-13'd134,  -13'd160,  13'd449,  -13'd251,  13'd449,  13'd652,  -13'd239,  -13'd349,  -13'd140,  -13'd106,  13'd416,  13'd113,  -13'd176,  13'd415,  13'd68,  -13'd269,  
-13'd142,  13'd387,  -13'd462,  -13'd960,  13'd599,  -13'd503,  -13'd814,  13'd84,  13'd53,  13'd34,  13'd82,  -13'd790,  13'd104,  13'd636,  13'd222,  -13'd490,  
-13'd535,  13'd305,  -13'd496,  -13'd202,  -13'd101,  13'd496,  -13'd75,  13'd54,  
-13'd31,  13'd358,  13'd538,  -13'd717,  -13'd290,  13'd160,  -13'd550,  -13'd719,  -13'd542,  13'd850,  -13'd279,  -13'd709,  13'd857,  13'd259,  13'd72,  -13'd393,  
-13'd25,  13'd564,  -13'd245,  13'd684,  13'd124,  13'd429,  -13'd55,  -13'd1291,  -13'd78,  13'd563,  13'd396,  -13'd777,  -13'd64,  -13'd470,  13'd45,  -13'd12,  
-13'd230,  13'd179,  13'd119,  13'd246,  -13'd469,  -13'd655,  -13'd641,  -13'd136,  13'd470,  -13'd158,  -13'd689,  -13'd21,  -13'd230,  13'd42,  13'd62,  -13'd20,  
13'd406,  -13'd490,  13'd171,  -13'd750,  13'd930,  13'd117,  -13'd994,  -13'd248,  13'd100,  13'd1115,  13'd356,  13'd40,  13'd890,  -13'd234,  -13'd598,  13'd242,  
-13'd570,  -13'd41,  -13'd161,  13'd470,  13'd448,  -13'd570,  -13'd254,  13'd557,  -13'd888,  -13'd526,  13'd1005,  13'd638,  13'd263,  -13'd622,  13'd443,  13'd666,  
13'd303,  -13'd482,  -13'd517,  13'd14,  13'd157,  13'd707,  13'd327,  -13'd288,  13'd242,  -13'd176,  -13'd459,  13'd221,  13'd262,  -13'd316,  -13'd750,  13'd635,  
13'd258,  -13'd67,  -13'd458,  -13'd650,  13'd911,  -13'd83,  13'd59,  13'd79,  -13'd464,  13'd828,  13'd488,  -13'd622,  -13'd266,  -13'd151,  -13'd321,  13'd301,  
13'd107,  -13'd462,  -13'd180,  -13'd243,  13'd784,  -13'd240,  13'd567,  13'd893,  
13'd557,  13'd153,  13'd894,  -13'd202,  13'd359,  13'd250,  13'd521,  -13'd877,  13'd78,  -13'd135,  -13'd121,  -13'd492,  13'd596,  -13'd131,  -13'd783,  13'd506,  
13'd183,  13'd525,  -13'd661,  -13'd359,  13'd290,  13'd11,  13'd535,  13'd801,  -13'd133,  13'd239,  -13'd267,  -13'd310,  -13'd232,  13'd311,  13'd172,  -13'd744,  
-13'd149,  -13'd267,  -13'd522,  -13'd615,  13'd792,  13'd322,  13'd438,  13'd279,  13'd214,  13'd226,  -13'd564,  -13'd636,  13'd243,  -13'd11,  13'd372,  13'd226,  
-13'd540,  -13'd718,  -13'd127,  -13'd263,  -13'd116,  13'd239,  13'd177,  13'd314,  -13'd1017,  13'd666,  13'd235,  -13'd294,  13'd625,  13'd259,  -13'd82,  13'd449,  
13'd656,  -13'd586,  13'd938,  13'd162,  -13'd61,  -13'd703,  13'd225,  -13'd257,  13'd494,  13'd246,  -13'd377,  -13'd559,  -13'd538,  -13'd32,  13'd176,  -13'd720,  
13'd108,  13'd441,  -13'd778,  -13'd122,  -13'd115,  -13'd49,  -13'd67,  13'd559,  13'd333,  13'd1059,  13'd295,  -13'd190,  -13'd240,  13'd336,  -13'd508,  -13'd2,  
-13'd26,  13'd133,  -13'd203,  -13'd86,  -13'd266,  13'd581,  13'd489,  13'd876,  -13'd333,  13'd636,  13'd11,  -13'd281,  -13'd230,  13'd110,  13'd20,  -13'd132,  
-13'd430,  -13'd1127,  13'd536,  13'd11,  13'd33,  -13'd69,  13'd37,  -13'd130,  
-13'd351,  13'd87,  13'd980,  -13'd16,  -13'd552,  -13'd97,  -13'd238,  -13'd393,  13'd68,  -13'd565,  13'd364,  -13'd1064,  -13'd414,  -13'd49,  -13'd491,  13'd281,  
-13'd171,  13'd900,  13'd605,  13'd106,  -13'd412,  -13'd561,  13'd93,  13'd1,  13'd709,  13'd138,  13'd833,  13'd99,  -13'd478,  13'd628,  -13'd490,  -13'd775,  
13'd805,  13'd60,  13'd576,  13'd533,  -13'd563,  -13'd133,  13'd116,  13'd290,  13'd383,  -13'd495,  -13'd718,  13'd531,  13'd553,  -13'd310,  -13'd5,  -13'd139,  
13'd657,  13'd13,  13'd239,  -13'd392,  -13'd304,  -13'd83,  -13'd496,  -13'd243,  -13'd659,  -13'd164,  13'd133,  13'd450,  13'd314,  13'd104,  -13'd432,  13'd447,  
-13'd62,  -13'd402,  -13'd192,  -13'd498,  13'd651,  13'd1107,  -13'd293,  13'd752,  -13'd593,  -13'd46,  13'd11,  -13'd221,  -13'd368,  -13'd355,  13'd146,  -13'd118,  
13'd478,  -13'd182,  -13'd297,  -13'd129,  13'd282,  -13'd173,  13'd417,  -13'd110,  13'd638,  -13'd429,  13'd66,  -13'd388,  13'd809,  13'd242,  13'd213,  13'd47,  
13'd331,  13'd160,  -13'd88,  13'd300,  -13'd289,  13'd131,  13'd75,  13'd933,  13'd227,  -13'd461,  13'd357,  -13'd604,  -13'd286,  13'd449,  13'd522,  13'd946,  
-13'd282,  -13'd215,  13'd727,  13'd654,  -13'd47,  -13'd341,  -13'd246,  13'd216,  
-13'd16,  13'd376,  13'd242,  -13'd286,  -13'd574,  13'd351,  13'd230,  13'd186,  13'd60,  13'd34,  -13'd81,  -13'd156,  -13'd501,  -13'd375,  -13'd101,  -13'd180,  
13'd323,  -13'd264,  13'd155,  -13'd248,  -13'd68,  -13'd592,  13'd51,  -13'd222,  13'd55,  -13'd630,  -13'd822,  13'd14,  13'd198,  13'd110,  -13'd345,  -13'd443,  
-13'd477,  13'd725,  13'd212,  -13'd364,  -13'd79,  -13'd508,  -13'd287,  -13'd273,  13'd323,  -13'd126,  -13'd88,  -13'd60,  13'd362,  -13'd416,  -13'd272,  13'd188,  
13'd146,  -13'd386,  -13'd237,  13'd262,  13'd165,  -13'd175,  -13'd207,  -13'd453,  -13'd164,  13'd320,  13'd134,  -13'd279,  13'd532,  -13'd534,  -13'd122,  -13'd637,  
-13'd444,  -13'd83,  13'd452,  13'd78,  13'd313,  -13'd46,  -13'd30,  -13'd45,  13'd252,  -13'd233,  13'd458,  13'd50,  -13'd124,  -13'd208,  -13'd162,  -13'd199,  
-13'd90,  -13'd136,  -13'd244,  13'd385,  13'd173,  -13'd637,  -13'd170,  -13'd264,  -13'd354,  13'd450,  -13'd670,  -13'd104,  -13'd306,  -13'd432,  13'd478,  -13'd29,  
13'd529,  13'd25,  13'd85,  13'd80,  -13'd451,  -13'd771,  -13'd71,  -13'd146,  -13'd644,  -13'd153,  -13'd159,  -13'd609,  -13'd165,  13'd45,  -13'd20,  13'd576,  
-13'd380,  -13'd96,  13'd85,  -13'd155,  -13'd450,  13'd206,  13'd30,  -13'd578,  
13'd16,  -13'd69,  -13'd151,  13'd479,  13'd110,  -13'd265,  -13'd642,  13'd230,  -13'd683,  -13'd325,  13'd2,  -13'd604,  -13'd181,  -13'd291,  13'd61,  13'd7,  
-13'd114,  -13'd424,  -13'd381,  13'd137,  -13'd140,  -13'd39,  -13'd62,  -13'd660,  -13'd38,  13'd259,  13'd403,  -13'd407,  13'd218,  -13'd419,  -13'd19,  13'd19,  
13'd181,  -13'd848,  -13'd62,  -13'd600,  -13'd594,  13'd65,  13'd327,  -13'd136,  -13'd529,  -13'd498,  13'd227,  -13'd18,  -13'd17,  -13'd291,  -13'd256,  -13'd37,  
13'd397,  13'd511,  -13'd297,  13'd619,  -13'd259,  -13'd767,  -13'd153,  -13'd45,  -13'd686,  13'd119,  13'd169,  -13'd808,  -13'd85,  -13'd316,  13'd700,  -13'd262,  
-13'd735,  -13'd571,  13'd303,  -13'd129,  -13'd257,  -13'd415,  13'd483,  -13'd348,  -13'd546,  -13'd144,  -13'd300,  -13'd68,  -13'd179,  -13'd815,  13'd173,  -13'd15,  
-13'd189,  -13'd92,  13'd280,  -13'd513,  -13'd408,  13'd303,  -13'd337,  -13'd683,  -13'd676,  -13'd681,  -13'd217,  -13'd297,  -13'd316,  13'd368,  13'd766,  -13'd18,  
13'd279,  -13'd339,  -13'd691,  -13'd51,  13'd549,  13'd406,  13'd535,  13'd215,  -13'd85,  13'd71,  -13'd93,  -13'd271,  13'd171,  13'd52,  -13'd852,  -13'd416,  
-13'd822,  -13'd764,  13'd198,  -13'd705,  -13'd337,  13'd155,  13'd149,  -13'd277,  
13'd18,  -13'd699,  -13'd590,  13'd385,  -13'd111,  13'd146,  -13'd124,  -13'd1602,  -13'd744,  -13'd358,  -13'd232,  13'd587,  -13'd81,  13'd203,  13'd426,  -13'd201,  
-13'd208,  -13'd128,  -13'd319,  -13'd147,  13'd141,  13'd217,  13'd483,  -13'd608,  -13'd297,  13'd931,  13'd767,  13'd618,  -13'd186,  13'd434,  13'd427,  13'd562,  
13'd258,  13'd883,  13'd534,  13'd313,  13'd336,  -13'd237,  13'd459,  -13'd413,  13'd459,  13'd724,  13'd53,  -13'd639,  -13'd870,  13'd382,  -13'd291,  -13'd865,  
13'd410,  -13'd416,  13'd148,  -13'd641,  13'd634,  13'd562,  13'd65,  -13'd21,  -13'd396,  13'd109,  13'd338,  13'd237,  13'd397,  -13'd113,  13'd406,  -13'd651,  
13'd170,  13'd416,  -13'd280,  -13'd1081,  -13'd112,  -13'd93,  13'd965,  -13'd324,  -13'd98,  -13'd432,  -13'd168,  -13'd550,  13'd207,  -13'd31,  -13'd476,  -13'd276,  
13'd581,  13'd172,  -13'd542,  -13'd616,  13'd530,  -13'd369,  -13'd708,  -13'd530,  -13'd294,  13'd1061,  13'd121,  13'd621,  13'd207,  -13'd357,  -13'd536,  13'd204,  
-13'd358,  -13'd294,  -13'd130,  -13'd109,  -13'd92,  -13'd893,  -13'd257,  -13'd573,  13'd262,  -13'd207,  13'd773,  -13'd267,  13'd137,  13'd1495,  -13'd48,  13'd528,  
-13'd352,  13'd271,  13'd1011,  -13'd77,  -13'd59,  13'd274,  13'd179,  13'd19,  
13'd495,  -13'd107,  13'd427,  13'd388,  -13'd120,  -13'd690,  -13'd125,  13'd58,  -13'd247,  13'd680,  13'd1119,  13'd451,  -13'd749,  -13'd607,  -13'd653,  13'd103,  
-13'd346,  -13'd273,  13'd502,  13'd7,  -13'd153,  -13'd474,  13'd563,  13'd464,  -13'd520,  13'd130,  13'd277,  13'd654,  -13'd813,  -13'd165,  13'd195,  13'd61,  
13'd61,  -13'd27,  13'd209,  13'd253,  13'd59,  13'd450,  13'd110,  13'd103,  -13'd106,  13'd196,  13'd358,  -13'd269,  -13'd791,  13'd26,  -13'd1412,  -13'd340,  
-13'd350,  13'd486,  -13'd7,  13'd846,  -13'd1054,  13'd223,  13'd752,  13'd503,  13'd643,  -13'd933,  -13'd540,  -13'd760,  13'd605,  -13'd492,  13'd411,  13'd260,  
13'd232,  -13'd170,  13'd171,  13'd722,  13'd155,  13'd341,  13'd586,  13'd284,  13'd91,  -13'd663,  -13'd557,  -13'd213,  -13'd806,  -13'd1177,  -13'd146,  -13'd172,  
13'd381,  13'd27,  -13'd304,  -13'd715,  13'd955,  13'd98,  13'd38,  -13'd171,  13'd332,  13'd42,  13'd823,  13'd333,  13'd54,  -13'd8,  -13'd628,  13'd61,  
13'd197,  -13'd178,  13'd935,  13'd1211,  -13'd330,  13'd1331,  -13'd120,  -13'd254,  13'd244,  -13'd220,  13'd250,  13'd236,  13'd157,  -13'd1001,  13'd399,  13'd309,  
13'd85,  -13'd428,  13'd286,  -13'd487,  -13'd163,  -13'd355,  13'd442,  -13'd259,  
-13'd73,  13'd293,  13'd174,  -13'd253,  13'd369,  -13'd352,  -13'd1,  13'd808,  13'd1208,  -13'd602,  13'd334,  -13'd520,  -13'd642,  -13'd820,  -13'd345,  -13'd100,  
13'd374,  -13'd158,  -13'd290,  13'd759,  -13'd67,  13'd222,  -13'd199,  -13'd170,  13'd15,  13'd225,  -13'd374,  -13'd437,  -13'd598,  13'd158,  13'd929,  13'd308,  
13'd133,  -13'd563,  -13'd311,  13'd304,  13'd1045,  13'd260,  13'd32,  13'd691,  13'd88,  13'd26,  13'd437,  -13'd621,  13'd269,  13'd280,  -13'd11,  13'd119,  
-13'd205,  13'd287,  13'd7,  -13'd243,  13'd396,  -13'd14,  13'd13,  13'd225,  13'd126,  -13'd598,  -13'd782,  -13'd297,  13'd470,  13'd179,  13'd372,  13'd190,  
-13'd470,  13'd288,  -13'd141,  -13'd10,  -13'd233,  13'd446,  -13'd134,  13'd106,  13'd832,  -13'd536,  -13'd599,  -13'd904,  -13'd55,  13'd645,  13'd393,  13'd765,  
13'd546,  13'd386,  -13'd346,  13'd1004,  -13'd78,  13'd193,  -13'd46,  13'd589,  13'd658,  13'd147,  -13'd462,  13'd491,  13'd756,  -13'd284,  -13'd135,  -13'd122,  
-13'd159,  13'd306,  -13'd1513,  -13'd646,  13'd265,  -13'd494,  -13'd988,  13'd1106,  13'd475,  -13'd495,  -13'd375,  -13'd464,  -13'd59,  -13'd660,  13'd132,  -13'd164,  
-13'd372,  13'd1136,  13'd483,  -13'd277,  -13'd246,  -13'd534,  13'd30,  13'd192,  
13'd64,  -13'd297,  -13'd956,  13'd282,  13'd560,  13'd217,  -13'd125,  -13'd500,  -13'd102,  13'd860,  -13'd1026,  13'd287,  13'd317,  13'd278,  13'd636,  -13'd499,  
13'd741,  13'd268,  13'd511,  13'd758,  13'd728,  13'd566,  13'd483,  13'd130,  13'd103,  -13'd788,  -13'd235,  13'd5,  13'd444,  -13'd299,  13'd763,  -13'd624,  
-13'd658,  -13'd595,  13'd487,  13'd122,  -13'd606,  -13'd200,  13'd129,  13'd300,  13'd866,  -13'd636,  -13'd235,  13'd199,  13'd211,  13'd665,  13'd643,  13'd835,  
13'd123,  -13'd631,  13'd499,  -13'd533,  13'd78,  -13'd28,  -13'd771,  13'd160,  13'd108,  13'd152,  -13'd1,  13'd305,  -13'd233,  13'd100,  -13'd820,  13'd358,  
-13'd522,  13'd216,  13'd172,  13'd234,  13'd452,  -13'd591,  -13'd193,  -13'd587,  -13'd534,  13'd467,  -13'd559,  13'd847,  13'd1058,  13'd635,  -13'd215,  -13'd53,  
-13'd278,  13'd91,  -13'd534,  -13'd468,  -13'd437,  13'd391,  13'd302,  13'd406,  13'd216,  -13'd259,  -13'd244,  13'd325,  13'd750,  13'd778,  13'd50,  -13'd168,  
13'd634,  -13'd797,  13'd428,  -13'd701,  -13'd6,  13'd189,  -13'd609,  -13'd714,  13'd152,  13'd56,  -13'd761,  13'd615,  -13'd215,  -13'd1109,  13'd322,  13'd550,  
-13'd323,  13'd222,  -13'd335,  13'd620,  13'd580,  13'd52,  -13'd402,  -13'd431,  
-13'd728,  -13'd208,  -13'd389,  -13'd27,  -13'd132,  -13'd341,  13'd697,  -13'd921,  13'd1126,  13'd345,  13'd468,  -13'd372,  -13'd159,  13'd540,  -13'd231,  13'd471,  
13'd342,  -13'd385,  13'd680,  13'd442,  13'd36,  13'd646,  13'd774,  -13'd785,  -13'd669,  -13'd253,  -13'd428,  -13'd507,  13'd838,  -13'd344,  -13'd574,  13'd981,  
13'd650,  -13'd25,  13'd180,  13'd374,  -13'd562,  13'd301,  13'd192,  -13'd216,  -13'd297,  13'd575,  13'd802,  13'd325,  -13'd192,  13'd180,  -13'd409,  -13'd62,  
-13'd414,  13'd148,  -13'd249,  13'd286,  -13'd87,  -13'd295,  13'd166,  13'd59,  13'd369,  -13'd209,  13'd87,  13'd1076,  -13'd178,  -13'd384,  13'd117,  13'd120,  
13'd6,  -13'd393,  -13'd70,  13'd589,  13'd403,  13'd1008,  -13'd320,  13'd522,  13'd544,  -13'd551,  13'd550,  -13'd723,  13'd307,  13'd151,  13'd628,  13'd680,  
-13'd517,  -13'd122,  13'd431,  13'd1168,  -13'd17,  -13'd254,  13'd493,  -13'd710,  13'd671,  -13'd1047,  -13'd678,  -13'd116,  13'd179,  13'd307,  13'd328,  -13'd282,  
13'd472,  13'd446,  -13'd837,  -13'd95,  -13'd349,  13'd151,  13'd41,  -13'd157,  13'd213,  13'd968,  -13'd76,  -13'd840,  13'd112,  13'd151,  -13'd528,  -13'd67,  
13'd301,  13'd655,  -13'd49,  -13'd293,  13'd77,  -13'd764,  13'd73,  -13'd645,  
13'd431,  13'd215,  13'd771,  13'd209,  -13'd264,  13'd153,  13'd514,  13'd1180,  -13'd86,  13'd644,  -13'd601,  -13'd220,  -13'd257,  -13'd59,  -13'd495,  -13'd931,  
-13'd756,  13'd434,  13'd233,  -13'd271,  -13'd347,  -13'd409,  -13'd357,  13'd456,  -13'd251,  -13'd189,  13'd599,  13'd62,  -13'd478,  13'd409,  -13'd191,  -13'd116,  
-13'd284,  -13'd95,  -13'd284,  13'd594,  13'd177,  13'd21,  13'd457,  13'd78,  13'd650,  -13'd149,  13'd163,  -13'd89,  13'd240,  -13'd222,  -13'd158,  13'd477,  
13'd456,  13'd776,  13'd31,  -13'd1122,  -13'd789,  -13'd384,  13'd247,  -13'd43,  13'd389,  -13'd159,  13'd802,  13'd109,  13'd223,  13'd286,  13'd493,  13'd419,  
-13'd594,  13'd221,  -13'd740,  -13'd761,  -13'd456,  -13'd458,  -13'd795,  13'd222,  -13'd749,  13'd150,  13'd410,  13'd17,  13'd902,  -13'd216,  13'd129,  13'd244,  
13'd473,  -13'd256,  13'd276,  13'd32,  13'd286,  13'd477,  13'd384,  13'd609,  13'd352,  -13'd207,  13'd653,  -13'd706,  -13'd79,  13'd674,  13'd252,  -13'd188,  
-13'd173,  -13'd91,  13'd431,  -13'd129,  13'd644,  13'd125,  13'd687,  13'd475,  13'd63,  -13'd355,  -13'd337,  -13'd770,  -13'd166,  -13'd1047,  -13'd280,  -13'd293,  
13'd272,  -13'd85,  -13'd411,  13'd195,  13'd159,  -13'd502,  13'd161,  13'd498,  
-13'd266,  13'd336,  13'd418,  -13'd95,  -13'd55,  -13'd234,  -13'd106,  13'd336,  -13'd59,  13'd830,  13'd415,  -13'd660,  13'd86,  -13'd454,  13'd226,  -13'd1337,  
-13'd132,  13'd524,  13'd65,  -13'd371,  13'd50,  -13'd41,  13'd270,  13'd384,  -13'd327,  -13'd184,  -13'd495,  -13'd1327,  -13'd36,  -13'd394,  13'd489,  13'd374,  
-13'd281,  13'd477,  -13'd278,  13'd387,  13'd74,  -13'd1465,  -13'd441,  -13'd348,  -13'd90,  -13'd642,  13'd490,  -13'd77,  13'd523,  13'd809,  -13'd28,  13'd322,  
13'd267,  13'd440,  13'd322,  -13'd304,  -13'd696,  -13'd692,  -13'd730,  13'd153,  -13'd207,  13'd621,  13'd423,  -13'd119,  -13'd880,  -13'd264,  -13'd537,  13'd47,  
13'd330,  13'd413,  -13'd33,  13'd331,  -13'd306,  13'd82,  13'd688,  -13'd195,  -13'd625,  -13'd810,  13'd193,  13'd385,  13'd451,  13'd694,  13'd40,  -13'd258,  
13'd107,  13'd132,  13'd617,  13'd580,  13'd211,  -13'd6,  -13'd926,  -13'd516,  13'd128,  -13'd618,  13'd340,  -13'd127,  -13'd61,  13'd637,  13'd31,  -13'd657,  
13'd845,  -13'd200,  13'd692,  -13'd307,  13'd27,  13'd22,  -13'd170,  13'd626,  13'd158,  13'd6,  -13'd428,  -13'd1330,  -13'd70,  -13'd316,  -13'd1129,  13'd608,  
-13'd357,  13'd615,  -13'd963,  -13'd219,  -13'd545,  -13'd302,  13'd430,  13'd395,  
-13'd36,  13'd509,  13'd201,  13'd28,  13'd455,  -13'd156,  -13'd224,  13'd1170,  13'd647,  -13'd264,  13'd18,  -13'd104,  13'd0,  13'd68,  13'd818,  13'd196,  
13'd39,  -13'd262,  -13'd335,  13'd694,  13'd702,  13'd198,  13'd532,  13'd83,  13'd323,  -13'd87,  -13'd84,  -13'd71,  13'd553,  13'd805,  13'd513,  13'd599,  
-13'd385,  -13'd147,  -13'd168,  13'd445,  -13'd691,  13'd414,  13'd29,  13'd727,  -13'd592,  -13'd280,  13'd811,  13'd230,  -13'd5,  13'd250,  13'd18,  13'd637,  
-13'd737,  13'd113,  -13'd9,  13'd582,  -13'd395,  13'd26,  -13'd384,  -13'd32,  13'd230,  -13'd1108,  -13'd168,  13'd570,  -13'd487,  13'd879,  13'd309,  13'd103,  
-13'd434,  -13'd276,  -13'd54,  13'd296,  13'd69,  -13'd111,  -13'd180,  -13'd267,  13'd330,  -13'd85,  -13'd25,  13'd29,  13'd297,  -13'd2,  -13'd185,  -13'd538,  
-13'd549,  13'd170,  13'd476,  13'd57,  -13'd78,  13'd133,  -13'd134,  -13'd261,  13'd390,  -13'd272,  13'd256,  13'd269,  -13'd13,  13'd6,  13'd225,  -13'd151,  
13'd188,  13'd523,  -13'd1310,  13'd238,  -13'd13,  -13'd343,  -13'd715,  -13'd474,  13'd31,  13'd277,  13'd38,  -13'd125,  -13'd239,  -13'd596,  -13'd756,  -13'd9,  
13'd501,  13'd1076,  -13'd189,  13'd164,  -13'd431,  13'd112,  13'd274,  -13'd587,  
-13'd405,  13'd293,  -13'd688,  13'd137,  -13'd57,  13'd128,  -13'd476,  -13'd1342,  -13'd1017,  -13'd636,  -13'd147,  -13'd601,  -13'd874,  -13'd84,  -13'd397,  -13'd50,  
-13'd513,  -13'd445,  -13'd38,  -13'd371,  -13'd492,  -13'd189,  -13'd58,  13'd198,  -13'd65,  -13'd408,  -13'd516,  -13'd52,  -13'd211,  -13'd436,  -13'd275,  -13'd12,  
-13'd119,  13'd592,  13'd487,  -13'd359,  13'd305,  -13'd180,  -13'd398,  13'd464,  -13'd350,  13'd53,  13'd129,  13'd474,  13'd260,  -13'd89,  -13'd278,  -13'd585,  
-13'd194,  -13'd127,  13'd279,  13'd312,  13'd144,  -13'd488,  13'd313,  -13'd355,  -13'd251,  -13'd774,  -13'd366,  -13'd669,  -13'd849,  -13'd269,  13'd36,  -13'd44,  
-13'd294,  13'd170,  13'd286,  13'd573,  13'd2,  -13'd194,  13'd923,  -13'd668,  13'd151,  -13'd415,  13'd498,  -13'd288,  -13'd402,  -13'd784,  -13'd738,  -13'd469,  
13'd6,  -13'd383,  13'd4,  -13'd494,  -13'd499,  -13'd521,  13'd330,  13'd147,  -13'd501,  -13'd220,  13'd242,  13'd223,  13'd183,  -13'd78,  13'd258,  -13'd392,  
-13'd826,  -13'd226,  13'd553,  13'd596,  13'd486,  -13'd43,  -13'd662,  -13'd920,  13'd76,  -13'd616,  -13'd287,  -13'd560,  13'd279,  -13'd261,  -13'd77,  -13'd549,  
-13'd21,  13'd130,  -13'd14,  13'd38,  -13'd185,  13'd61,  -13'd0,  -13'd601,  
-13'd30,  13'd481,  13'd178,  -13'd476,  13'd33,  -13'd359,  13'd219,  -13'd175,  13'd124,  13'd27,  13'd497,  -13'd353,  -13'd431,  -13'd359,  -13'd118,  -13'd10,  
13'd912,  13'd343,  -13'd32,  13'd667,  -13'd289,  13'd396,  -13'd117,  -13'd1446,  13'd121,  -13'd333,  13'd352,  13'd539,  -13'd122,  -13'd95,  13'd589,  -13'd441,  
13'd142,  13'd267,  -13'd525,  13'd530,  -13'd497,  13'd493,  -13'd93,  13'd78,  -13'd814,  13'd584,  -13'd74,  13'd415,  -13'd589,  13'd676,  13'd33,  13'd72,  
13'd284,  13'd673,  13'd698,  -13'd164,  -13'd91,  13'd114,  13'd875,  -13'd449,  13'd491,  -13'd622,  -13'd378,  -13'd971,  13'd109,  13'd197,  13'd235,  -13'd652,  
-13'd481,  13'd696,  13'd135,  13'd213,  -13'd110,  -13'd755,  13'd194,  13'd234,  13'd850,  -13'd348,  13'd149,  -13'd470,  -13'd1080,  -13'd150,  -13'd844,  -13'd206,  
13'd298,  -13'd20,  13'd273,  -13'd109,  13'd932,  13'd686,  13'd293,  -13'd296,  -13'd531,  -13'd832,  13'd7,  13'd500,  -13'd360,  13'd140,  13'd47,  -13'd346,  
13'd207,  -13'd138,  -13'd292,  13'd19,  13'd733,  13'd289,  -13'd445,  -13'd407,  13'd746,  -13'd330,  13'd70,  13'd299,  -13'd299,  13'd1275,  -13'd398,  -13'd372,  
13'd122,  13'd649,  -13'd15,  -13'd682,  -13'd372,  13'd442,  13'd131,  -13'd31,  
-13'd715,  13'd44,  -13'd617,  13'd326,  13'd226,  13'd580,  13'd91,  13'd488,  -13'd830,  13'd742,  -13'd1018,  13'd383,  13'd148,  13'd729,  13'd366,  -13'd857,  
13'd743,  13'd665,  -13'd252,  -13'd417,  -13'd378,  13'd123,  13'd317,  13'd399,  -13'd137,  -13'd6,  -13'd184,  13'd293,  13'd1114,  13'd476,  13'd1336,  13'd139,  
-13'd219,  13'd711,  13'd183,  13'd196,  13'd114,  -13'd575,  -13'd96,  -13'd80,  13'd278,  -13'd446,  -13'd656,  -13'd633,  -13'd106,  13'd144,  -13'd266,  13'd343,  
-13'd643,  -13'd174,  -13'd20,  -13'd163,  13'd192,  -13'd565,  -13'd1114,  13'd321,  13'd131,  13'd681,  13'd225,  13'd273,  -13'd225,  13'd343,  -13'd73,  -13'd116,  
-13'd180,  13'd322,  -13'd452,  -13'd363,  -13'd28,  -13'd567,  -13'd119,  13'd343,  -13'd417,  -13'd145,  -13'd84,  13'd379,  -13'd224,  13'd431,  -13'd526,  13'd322,  
13'd381,  13'd302,  13'd355,  13'd406,  -13'd163,  -13'd476,  -13'd100,  13'd410,  13'd327,  -13'd398,  -13'd912,  13'd702,  -13'd587,  -13'd0,  13'd767,  13'd148,  
13'd391,  -13'd349,  13'd35,  -13'd377,  13'd374,  13'd24,  -13'd505,  -13'd857,  -13'd73,  13'd184,  13'd116,  13'd284,  -13'd229,  -13'd422,  13'd157,  -13'd551,  
13'd1066,  -13'd269,  -13'd589,  13'd20,  13'd436,  -13'd512,  13'd116,  -13'd450,  
13'd618,  -13'd23,  13'd704,  13'd103,  -13'd373,  13'd664,  -13'd700,  13'd422,  -13'd547,  -13'd652,  13'd98,  13'd154,  -13'd439,  13'd86,  13'd215,  -13'd123,  
13'd422,  -13'd360,  13'd391,  13'd395,  -13'd376,  -13'd311,  13'd94,  -13'd31,  -13'd123,  -13'd44,  13'd746,  13'd614,  -13'd779,  -13'd178,  -13'd11,  13'd6,  
-13'd129,  -13'd306,  13'd36,  13'd466,  13'd567,  -13'd407,  13'd127,  -13'd616,  13'd627,  13'd811,  13'd929,  -13'd273,  -13'd151,  -13'd635,  13'd139,  -13'd514,  
13'd31,  13'd116,  13'd244,  13'd527,  13'd115,  -13'd48,  13'd298,  -13'd712,  -13'd709,  13'd35,  -13'd387,  -13'd786,  13'd103,  -13'd258,  13'd553,  13'd48,  
13'd83,  13'd678,  13'd254,  -13'd34,  13'd383,  13'd789,  13'd288,  13'd65,  13'd529,  -13'd269,  -13'd236,  13'd174,  -13'd122,  -13'd693,  -13'd987,  -13'd629,  
-13'd334,  13'd344,  -13'd142,  -13'd553,  13'd581,  13'd265,  13'd354,  13'd30,  13'd563,  13'd878,  13'd284,  13'd199,  -13'd301,  13'd758,  -13'd137,  13'd896,  
-13'd242,  -13'd734,  13'd296,  -13'd124,  13'd207,  -13'd466,  13'd178,  13'd1033,  13'd189,  -13'd13,  -13'd202,  13'd856,  13'd557,  13'd471,  13'd1038,  13'd198,  
-13'd192,  -13'd70,  13'd866,  13'd27,  13'd43,  -13'd652,  -13'd844,  13'd358,  
-13'd794,  13'd370,  -13'd37,  -13'd356,  -13'd335,  13'd655,  13'd312,  -13'd222,  13'd161,  -13'd170,  -13'd569,  -13'd254,  -13'd503,  13'd158,  -13'd234,  13'd18,  
-13'd72,  13'd633,  13'd360,  13'd116,  13'd579,  -13'd605,  -13'd301,  13'd450,  -13'd430,  13'd168,  -13'd202,  -13'd629,  -13'd582,  -13'd75,  13'd38,  13'd482,  
-13'd340,  13'd229,  13'd71,  13'd0,  -13'd102,  -13'd588,  -13'd54,  -13'd425,  13'd186,  13'd40,  -13'd107,  -13'd116,  -13'd188,  -13'd111,  13'd248,  -13'd301,  
13'd111,  -13'd438,  13'd741,  -13'd160,  -13'd235,  -13'd777,  13'd244,  13'd314,  -13'd124,  -13'd399,  13'd422,  -13'd876,  -13'd93,  -13'd103,  -13'd368,  13'd83,  
13'd133,  -13'd184,  -13'd75,  -13'd260,  13'd223,  13'd91,  13'd183,  13'd406,  -13'd64,  13'd530,  -13'd16,  -13'd584,  -13'd142,  -13'd44,  -13'd554,  13'd353,  
13'd148,  -13'd268,  -13'd430,  -13'd221,  -13'd185,  -13'd192,  -13'd165,  13'd159,  13'd2,  -13'd174,  -13'd336,  -13'd479,  -13'd329,  -13'd411,  -13'd25,  13'd54,  
13'd208,  -13'd492,  -13'd703,  13'd503,  -13'd343,  -13'd337,  -13'd345,  -13'd804,  -13'd89,  13'd55,  -13'd91,  -13'd277,  -13'd76,  -13'd173,  -13'd344,  13'd665,  
13'd278,  13'd449,  13'd447,  13'd215,  -13'd360,  13'd122,  13'd216,  -13'd395,  
13'd833,  13'd275,  -13'd778,  -13'd348,  13'd67,  -13'd446,  -13'd28,  13'd358,  -13'd222,  -13'd550,  -13'd1125,  -13'd455,  13'd517,  -13'd394,  13'd354,  -13'd4,  
13'd821,  -13'd142,  13'd161,  13'd1056,  -13'd628,  13'd358,  13'd777,  13'd1157,  13'd31,  -13'd286,  13'd158,  -13'd332,  13'd97,  13'd56,  13'd814,  -13'd75,  
13'd34,  -13'd433,  -13'd510,  13'd497,  -13'd438,  13'd717,  13'd943,  -13'd330,  13'd437,  13'd10,  13'd283,  13'd117,  -13'd475,  -13'd643,  -13'd206,  13'd125,  
13'd173,  -13'd32,  -13'd409,  13'd537,  13'd359,  -13'd632,  -13'd104,  13'd55,  13'd85,  13'd472,  -13'd441,  -13'd764,  -13'd447,  -13'd168,  -13'd869,  13'd124,  
13'd714,  -13'd260,  13'd311,  13'd1186,  -13'd725,  13'd178,  -13'd123,  13'd307,  13'd192,  -13'd116,  -13'd330,  -13'd387,  13'd43,  -13'd85,  13'd282,  13'd47,  
-13'd92,  13'd594,  -13'd108,  13'd411,  13'd343,  -13'd277,  13'd597,  -13'd161,  13'd748,  13'd565,  -13'd167,  13'd96,  13'd212,  13'd650,  -13'd491,  13'd411,  
13'd412,  -13'd383,  -13'd2,  13'd824,  13'd122,  -13'd28,  13'd337,  13'd931,  -13'd118,  13'd11,  13'd504,  13'd283,  13'd727,  13'd506,  13'd844,  13'd68,  
-13'd67,  13'd528,  13'd254,  13'd505,  13'd688,  13'd653,  13'd335,  13'd48,  
13'd270,  13'd359,  -13'd829,  13'd337,  13'd227,  13'd389,  13'd33,  13'd404,  13'd276,  13'd137,  -13'd759,  -13'd479,  13'd625,  -13'd744,  13'd46,  13'd442,  
13'd527,  -13'd361,  13'd73,  -13'd576,  13'd147,  13'd55,  13'd641,  13'd472,  13'd675,  -13'd446,  -13'd272,  13'd162,  13'd470,  -13'd196,  13'd418,  13'd263,  
13'd252,  13'd446,  13'd523,  -13'd66,  -13'd762,  -13'd369,  -13'd111,  13'd215,  -13'd115,  -13'd267,  13'd187,  -13'd484,  13'd941,  13'd442,  -13'd300,  -13'd184,  
13'd252,  -13'd74,  13'd307,  -13'd142,  -13'd584,  -13'd548,  -13'd291,  -13'd389,  13'd989,  -13'd259,  -13'd578,  13'd192,  -13'd4,  13'd533,  -13'd218,  13'd11,  
-13'd636,  13'd1102,  13'd340,  -13'd112,  13'd53,  -13'd582,  13'd306,  -13'd660,  13'd271,  13'd31,  13'd670,  13'd177,  13'd758,  -13'd12,  13'd592,  -13'd176,  
13'd22,  13'd851,  13'd146,  13'd153,  -13'd747,  -13'd289,  13'd317,  -13'd275,  -13'd429,  -13'd344,  -13'd24,  -13'd154,  -13'd146,  -13'd97,  -13'd189,  13'd486,  
-13'd58,  13'd259,  -13'd5,  -13'd332,  13'd483,  13'd257,  13'd335,  -13'd722,  -13'd651,  13'd531,  13'd895,  -13'd1048,  13'd402,  13'd293,  -13'd56,  13'd443,  
-13'd214,  -13'd340,  -13'd27,  13'd452,  -13'd199,  -13'd798,  -13'd89,  13'd51,  
13'd201,  -13'd236,  13'd39,  13'd234,  -13'd569,  -13'd284,  -13'd122,  -13'd255,  13'd30,  -13'd114,  -13'd890,  13'd870,  13'd780,  13'd346,  13'd439,  13'd380,  
-13'd34,  13'd535,  -13'd15,  -13'd205,  13'd146,  -13'd316,  13'd529,  13'd424,  -13'd360,  13'd191,  -13'd124,  -13'd374,  13'd375,  13'd340,  -13'd650,  13'd885,  
13'd88,  13'd186,  13'd200,  13'd465,  13'd813,  -13'd662,  -13'd253,  13'd139,  13'd786,  13'd429,  -13'd538,  13'd236,  -13'd926,  -13'd142,  13'd82,  -13'd948,  
13'd212,  -13'd934,  13'd412,  13'd995,  -13'd785,  13'd629,  13'd552,  -13'd291,  13'd59,  13'd85,  -13'd380,  -13'd384,  13'd310,  -13'd272,  -13'd603,  -13'd408,  
-13'd184,  -13'd43,  13'd406,  -13'd87,  -13'd134,  -13'd549,  -13'd266,  13'd567,  13'd222,  13'd251,  13'd535,  13'd152,  13'd518,  -13'd151,  13'd575,  13'd158,  
-13'd273,  -13'd747,  -13'd35,  -13'd845,  -13'd219,  13'd395,  13'd592,  13'd427,  13'd599,  -13'd8,  13'd388,  13'd402,  -13'd673,  13'd745,  13'd80,  -13'd121,  
13'd127,  -13'd159,  13'd497,  -13'd605,  -13'd145,  -13'd43,  -13'd18,  -13'd572,  13'd469,  13'd84,  13'd1227,  13'd64,  -13'd95,  13'd875,  -13'd357,  13'd980,  
13'd799,  -13'd526,  13'd427,  13'd542,  13'd232,  -13'd379,  -13'd224,  -13'd141,  
13'd124,  13'd158,  13'd665,  13'd113,  13'd305,  13'd104,  13'd637,  13'd119,  13'd143,  -13'd87,  13'd331,  -13'd46,  13'd158,  13'd69,  -13'd477,  -13'd20,  
13'd166,  13'd270,  13'd616,  13'd330,  13'd486,  13'd153,  -13'd507,  -13'd716,  13'd174,  13'd10,  -13'd425,  13'd81,  13'd220,  13'd5,  -13'd561,  -13'd320,  
13'd189,  13'd717,  -13'd228,  -13'd401,  13'd501,  -13'd91,  -13'd574,  -13'd430,  -13'd247,  -13'd269,  13'd1201,  13'd885,  -13'd104,  13'd230,  13'd205,  -13'd454,  
-13'd54,  13'd859,  13'd250,  13'd653,  -13'd571,  13'd437,  -13'd551,  -13'd104,  13'd60,  -13'd2,  -13'd583,  -13'd356,  13'd491,  -13'd219,  13'd1030,  -13'd826,  
-13'd773,  13'd335,  13'd362,  -13'd277,  13'd189,  13'd234,  -13'd143,  -13'd32,  13'd791,  -13'd386,  -13'd4,  13'd858,  -13'd37,  13'd421,  -13'd57,  -13'd527,  
13'd11,  -13'd144,  13'd1054,  13'd727,  13'd146,  13'd97,  13'd207,  -13'd641,  -13'd6,  13'd196,  13'd167,  -13'd279,  -13'd363,  13'd598,  -13'd227,  -13'd307,  
13'd239,  -13'd475,  13'd744,  13'd519,  13'd710,  13'd681,  -13'd129,  -13'd124,  -13'd440,  13'd529,  -13'd356,  -13'd342,  -13'd28,  -13'd218,  -13'd662,  13'd923,  
13'd207,  -13'd47,  13'd460,  -13'd172,  -13'd192,  -13'd184,  -13'd291,  -13'd88,  
13'd429,  -13'd16,  -13'd821,  13'd280,  -13'd586,  -13'd214,  13'd463,  -13'd9,  13'd475,  13'd761,  13'd313,  13'd264,  -13'd162,  13'd946,  13'd137,  -13'd1270,  
-13'd1026,  -13'd33,  -13'd776,  13'd759,  13'd135,  13'd48,  13'd322,  -13'd503,  13'd343,  -13'd161,  13'd933,  -13'd103,  13'd97,  13'd1154,  13'd248,  13'd383,  
-13'd352,  -13'd647,  -13'd755,  -13'd700,  13'd514,  -13'd217,  -13'd28,  -13'd150,  13'd472,  13'd205,  -13'd826,  -13'd607,  13'd194,  13'd627,  -13'd521,  13'd807,  
13'd67,  -13'd938,  -13'd95,  -13'd308,  -13'd15,  -13'd674,  -13'd79,  -13'd69,  13'd226,  13'd1097,  13'd44,  -13'd262,  13'd532,  13'd128,  -13'd448,  -13'd688,  
13'd633,  -13'd250,  13'd430,  13'd483,  -13'd233,  -13'd219,  -13'd975,  13'd106,  -13'd109,  13'd334,  -13'd259,  13'd774,  13'd645,  -13'd134,  13'd205,  -13'd417,  
-13'd278,  -13'd323,  -13'd135,  13'd459,  13'd97,  13'd60,  -13'd945,  13'd357,  -13'd235,  13'd440,  -13'd457,  13'd566,  13'd351,  -13'd177,  -13'd502,  -13'd527,  
-13'd248,  -13'd287,  -13'd73,  -13'd751,  13'd457,  -13'd1237,  13'd652,  13'd1226,  13'd274,  -13'd79,  -13'd529,  13'd215,  13'd82,  13'd536,  13'd714,  -13'd583,  
-13'd381,  13'd579,  13'd760,  13'd304,  13'd60,  -13'd733,  -13'd480,  -13'd391,  
13'd25,  13'd109,  -13'd383,  13'd112,  13'd372,  -13'd90,  -13'd977,  -13'd419,  13'd299,  -13'd15,  13'd324,  -13'd197,  -13'd250,  -13'd151,  -13'd195,  -13'd609,  
-13'd757,  13'd371,  -13'd221,  13'd39,  -13'd398,  -13'd276,  13'd65,  13'd237,  13'd234,  -13'd397,  13'd43,  -13'd221,  13'd32,  -13'd211,  -13'd35,  -13'd538,  
13'd326,  -13'd725,  13'd457,  13'd13,  -13'd44,  -13'd583,  13'd86,  -13'd942,  13'd102,  -13'd60,  13'd637,  -13'd674,  -13'd884,  13'd349,  -13'd225,  -13'd155,  
-13'd378,  13'd261,  13'd31,  -13'd452,  -13'd23,  -13'd521,  -13'd356,  -13'd191,  -13'd343,  13'd105,  -13'd741,  -13'd657,  -13'd323,  -13'd718,  -13'd109,  -13'd561,  
-13'd42,  -13'd344,  13'd66,  -13'd744,  13'd33,  -13'd295,  -13'd947,  -13'd404,  -13'd103,  -13'd714,  -13'd249,  -13'd242,  13'd375,  13'd327,  -13'd4,  13'd364,  
-13'd687,  -13'd328,  -13'd953,  -13'd7,  -13'd665,  -13'd464,  -13'd995,  -13'd179,  -13'd85,  13'd58,  -13'd6,  -13'd113,  -13'd497,  -13'd653,  -13'd137,  13'd415,  
-13'd548,  -13'd443,  -13'd308,  13'd20,  -13'd832,  13'd74,  13'd556,  -13'd309,  13'd100,  -13'd541,  -13'd13,  -13'd266,  -13'd553,  -13'd540,  -13'd223,  -13'd150,  
-13'd240,  13'd166,  -13'd45,  -13'd104,  13'd177,  13'd139,  -13'd306,  13'd448,  
13'd1185,  -13'd129,  13'd711,  -13'd200,  13'd1015,  -13'd179,  -13'd238,  13'd329,  -13'd990,  -13'd114,  -13'd166,  13'd257,  -13'd816,  13'd924,  -13'd78,  -13'd616,  
13'd977,  13'd191,  -13'd84,  13'd169,  13'd130,  -13'd257,  -13'd499,  13'd388,  13'd18,  13'd895,  13'd176,  -13'd781,  -13'd515,  13'd557,  -13'd112,  13'd416,  
-13'd121,  13'd110,  13'd80,  -13'd290,  -13'd20,  13'd615,  13'd140,  13'd126,  13'd534,  13'd336,  13'd884,  -13'd234,  13'd80,  13'd101,  13'd27,  -13'd898,  
13'd279,  -13'd116,  13'd786,  13'd865,  -13'd1,  13'd802,  13'd238,  -13'd57,  13'd35,  -13'd157,  -13'd151,  -13'd73,  13'd491,  13'd118,  -13'd576,  -13'd968,  
13'd132,  -13'd190,  -13'd147,  -13'd836,  -13'd262,  13'd118,  13'd328,  13'd389,  13'd571,  13'd205,  13'd565,  -13'd426,  13'd241,  13'd462,  13'd676,  13'd330,  
-13'd444,  13'd440,  13'd19,  -13'd12,  -13'd55,  -13'd433,  -13'd709,  -13'd381,  -13'd714,  -13'd51,  13'd890,  -13'd28,  -13'd202,  13'd150,  13'd376,  -13'd941,  
-13'd504,  -13'd583,  13'd113,  13'd372,  13'd687,  13'd598,  13'd196,  -13'd116,  13'd370,  13'd191,  13'd309,  13'd21,  13'd604,  -13'd1018,  13'd27,  13'd398,  
-13'd302,  13'd932,  -13'd428,  13'd525,  13'd20,  -13'd222,  -13'd229,  13'd130,  
-13'd514,  -13'd320,  -13'd4,  -13'd460,  13'd193,  -13'd264,  13'd421,  13'd34,  13'd325,  -13'd302,  -13'd469,  13'd93,  -13'd63,  -13'd80,  -13'd298,  13'd1,  
-13'd423,  13'd302,  13'd459,  -13'd520,  -13'd339,  13'd257,  -13'd189,  13'd553,  -13'd197,  13'd443,  13'd642,  13'd257,  -13'd86,  13'd527,  -13'd429,  -13'd475,  
13'd115,  -13'd195,  13'd196,  -13'd145,  -13'd331,  13'd448,  13'd644,  -13'd142,  -13'd227,  13'd225,  -13'd474,  13'd710,  -13'd52,  -13'd397,  -13'd71,  13'd664,  
13'd229,  13'd72,  -13'd300,  -13'd1087,  13'd82,  -13'd122,  -13'd129,  13'd77,  13'd612,  -13'd621,  -13'd740,  -13'd627,  13'd367,  -13'd104,  -13'd1140,  13'd101,  
13'd324,  -13'd709,  13'd3,  13'd696,  13'd786,  13'd52,  13'd53,  13'd505,  13'd379,  13'd127,  13'd90,  13'd473,  -13'd935,  -13'd56,  13'd402,  -13'd396,  
13'd610,  13'd22,  -13'd9,  13'd509,  13'd91,  -13'd756,  13'd388,  13'd705,  -13'd270,  13'd357,  13'd901,  13'd331,  -13'd44,  13'd13,  -13'd307,  13'd429,  
-13'd359,  -13'd84,  -13'd180,  13'd181,  -13'd301,  13'd387,  -13'd359,  13'd1260,  13'd69,  13'd431,  -13'd138,  -13'd370,  13'd204,  -13'd675,  -13'd61,  13'd348,  
-13'd499,  13'd166,  -13'd603,  -13'd437,  13'd117,  13'd549,  13'd19,  13'd368,  
-13'd28,  13'd31,  -13'd555,  -13'd750,  13'd546,  13'd987,  13'd51,  -13'd468,  -13'd258,  -13'd628,  13'd136,  13'd304,  13'd313,  13'd695,  13'd272,  13'd572,  
13'd404,  13'd61,  -13'd766,  -13'd767,  13'd129,  -13'd138,  -13'd403,  13'd378,  13'd570,  -13'd867,  -13'd24,  -13'd528,  -13'd396,  13'd475,  13'd259,  13'd42,  
-13'd231,  13'd243,  -13'd409,  13'd67,  13'd35,  13'd188,  -13'd570,  13'd186,  -13'd469,  13'd624,  -13'd197,  -13'd69,  -13'd147,  13'd173,  -13'd293,  -13'd642,  
13'd434,  13'd260,  13'd198,  -13'd1150,  -13'd4,  -13'd357,  13'd455,  -13'd257,  -13'd46,  -13'd61,  -13'd464,  -13'd483,  -13'd677,  13'd330,  -13'd248,  13'd297,  
13'd588,  -13'd19,  -13'd359,  13'd84,  13'd252,  -13'd1285,  13'd518,  13'd236,  13'd675,  -13'd990,  13'd428,  -13'd121,  13'd111,  -13'd170,  13'd115,  -13'd592,  
13'd40,  13'd258,  13'd449,  -13'd681,  13'd316,  13'd449,  13'd173,  -13'd158,  13'd763,  13'd150,  13'd324,  13'd338,  13'd318,  -13'd263,  -13'd346,  13'd147,  
-13'd172,  -13'd17,  13'd710,  13'd659,  13'd394,  13'd102,  -13'd167,  -13'd344,  -13'd76,  13'd487,  13'd721,  -13'd211,  -13'd499,  -13'd213,  13'd63,  -13'd90,  
13'd32,  13'd80,  -13'd244,  -13'd86,  -13'd267,  -13'd441,  13'd136,  13'd567,  
13'd11,  -13'd15,  13'd43,  -13'd138,  13'd364,  -13'd232,  -13'd945,  13'd566,  -13'd1233,  -13'd154,  -13'd760,  -13'd390,  13'd267,  13'd463,  13'd358,  13'd42,  
-13'd486,  13'd731,  -13'd875,  -13'd174,  -13'd547,  -13'd486,  13'd180,  13'd992,  -13'd15,  13'd505,  -13'd70,  -13'd877,  13'd456,  13'd686,  -13'd686,  13'd966,  
-13'd771,  -13'd8,  13'd255,  13'd300,  13'd1121,  13'd537,  13'd117,  -13'd281,  13'd228,  13'd123,  -13'd172,  -13'd578,  13'd35,  -13'd692,  -13'd447,  -13'd1253,  
13'd431,  -13'd362,  -13'd755,  13'd230,  13'd391,  13'd84,  -13'd810,  13'd10,  -13'd366,  -13'd193,  13'd417,  13'd97,  -13'd166,  13'd535,  -13'd392,  13'd26,  
13'd592,  -13'd192,  -13'd264,  13'd133,  -13'd77,  -13'd593,  13'd300,  -13'd111,  13'd206,  -13'd494,  13'd367,  -13'd111,  -13'd1054,  13'd282,  13'd93,  -13'd439,  
-13'd390,  13'd316,  -13'd966,  -13'd39,  -13'd353,  13'd25,  -13'd306,  -13'd275,  -13'd27,  -13'd93,  -13'd103,  -13'd342,  -13'd75,  -13'd460,  -13'd385,  13'd385,  
13'd211,  -13'd314,  -13'd212,  -13'd1224,  13'd46,  -13'd13,  -13'd54,  13'd15,  -13'd335,  13'd519,  13'd98,  -13'd915,  -13'd335,  13'd865,  13'd211,  13'd809,  
-13'd383,  -13'd531,  13'd425,  13'd106,  13'd216,  13'd160,  13'd896,  13'd194,  
-13'd394,  -13'd633,  -13'd310,  -13'd201,  13'd278,  13'd21,  13'd76,  13'd34,  -13'd74,  13'd690,  -13'd262,  13'd584,  13'd74,  13'd172,  -13'd502,  13'd166,  
-13'd40,  -13'd64,  13'd6,  -13'd50,  -13'd313,  -13'd435,  -13'd474,  13'd403,  -13'd250,  13'd69,  13'd154,  13'd553,  -13'd81,  -13'd345,  -13'd683,  13'd435,  
-13'd913,  -13'd1,  13'd547,  -13'd96,  -13'd709,  -13'd128,  13'd351,  13'd426,  13'd450,  -13'd496,  13'd709,  13'd702,  -13'd238,  -13'd114,  -13'd421,  13'd271,  
13'd22,  13'd27,  13'd229,  13'd14,  13'd229,  -13'd362,  -13'd111,  -13'd276,  -13'd450,  13'd397,  13'd660,  13'd48,  13'd548,  -13'd246,  13'd69,  -13'd698,  
-13'd117,  13'd80,  13'd174,  13'd30,  13'd211,  -13'd220,  -13'd222,  13'd9,  -13'd304,  13'd1247,  13'd5,  13'd55,  13'd51,  -13'd18,  -13'd701,  13'd518,  
13'd7,  -13'd284,  -13'd571,  -13'd451,  -13'd273,  -13'd76,  -13'd765,  13'd678,  -13'd73,  13'd400,  13'd841,  13'd582,  13'd318,  13'd397,  -13'd510,  13'd716,  
-13'd583,  -13'd265,  13'd998,  13'd224,  13'd197,  13'd373,  13'd323,  13'd293,  -13'd800,  -13'd40,  -13'd19,  13'd916,  13'd40,  13'd185,  13'd186,  13'd170,  
13'd244,  -13'd528,  -13'd420,  13'd51,  13'd767,  13'd893,  -13'd177,  -13'd14,  
-13'd587,  -13'd303,  -13'd220,  -13'd116,  13'd687,  -13'd330,  13'd580,  13'd489,  13'd1124,  -13'd289,  13'd442,  -13'd217,  13'd127,  13'd378,  13'd853,  13'd208,  
13'd49,  -13'd470,  -13'd23,  -13'd305,  -13'd51,  -13'd136,  13'd286,  13'd421,  -13'd114,  13'd1084,  13'd77,  13'd526,  13'd0,  13'd94,  -13'd312,  -13'd712,  
13'd913,  -13'd125,  13'd276,  13'd163,  -13'd680,  13'd83,  -13'd228,  13'd95,  -13'd510,  -13'd193,  13'd490,  13'd19,  13'd1043,  13'd240,  -13'd599,  13'd439,  
13'd32,  13'd219,  13'd49,  13'd286,  -13'd673,  13'd577,  -13'd1098,  -13'd113,  13'd196,  -13'd936,  13'd243,  -13'd74,  -13'd274,  13'd452,  13'd804,  13'd874,  
13'd282,  13'd375,  13'd252,  -13'd306,  13'd565,  13'd159,  13'd451,  13'd45,  13'd436,  13'd308,  13'd41,  13'd157,  13'd359,  -13'd84,  -13'd424,  13'd77,  
-13'd681,  -13'd29,  13'd668,  13'd973,  13'd330,  13'd626,  13'd0,  -13'd543,  -13'd343,  13'd177,  13'd537,  -13'd258,  13'd742,  13'd323,  -13'd251,  -13'd519,  
-13'd299,  -13'd431,  -13'd313,  13'd1123,  -13'd489,  13'd572,  13'd312,  -13'd222,  13'd489,  -13'd448,  -13'd177,  13'd488,  -13'd20,  -13'd583,  -13'd357,  -13'd97,  
13'd392,  13'd894,  -13'd963,  13'd125,  -13'd299,  -13'd505,  13'd231,  -13'd510,  
-13'd22,  -13'd120,  -13'd795,  13'd359,  -13'd251,  13'd315,  13'd326,  -13'd2,  -13'd50,  13'd120,  -13'd209,  13'd42,  -13'd104,  13'd41,  13'd404,  -13'd325,  
-13'd708,  -13'd247,  13'd769,  13'd132,  13'd60,  -13'd376,  -13'd162,  -13'd601,  -13'd583,  -13'd22,  13'd639,  13'd391,  -13'd420,  13'd256,  -13'd282,  -13'd373,  
-13'd996,  13'd763,  -13'd332,  13'd76,  -13'd6,  13'd71,  -13'd239,  13'd72,  13'd615,  -13'd518,  -13'd517,  13'd164,  13'd38,  13'd246,  13'd825,  13'd897,  
13'd603,  -13'd500,  13'd905,  -13'd75,  13'd176,  13'd623,  -13'd197,  13'd3,  -13'd104,  13'd668,  13'd590,  13'd164,  13'd392,  -13'd8,  13'd1309,  13'd54,  
-13'd452,  -13'd104,  13'd198,  -13'd58,  13'd191,  -13'd164,  13'd354,  -13'd70,  13'd69,  13'd92,  -13'd733,  13'd693,  13'd179,  -13'd800,  -13'd369,  -13'd414,  
13'd165,  -13'd223,  13'd452,  -13'd460,  -13'd718,  13'd565,  -13'd302,  -13'd266,  13'd388,  13'd877,  13'd192,  13'd682,  -13'd516,  13'd55,  13'd252,  13'd708,  
-13'd47,  -13'd506,  13'd1112,  -13'd383,  13'd215,  -13'd156,  -13'd71,  13'd811,  -13'd629,  -13'd192,  -13'd242,  13'd309,  13'd291,  13'd239,  13'd436,  -13'd207,  
13'd147,  -13'd239,  13'd852,  -13'd44,  -13'd37,  13'd166,  13'd63,  -13'd76,  
13'd304,  -13'd563,  13'd402,  -13'd229,  13'd222,  13'd70,  -13'd211,  -13'd58,  13'd252,  13'd59,  -13'd598,  -13'd1,  13'd663,  13'd19,  13'd764,  -13'd38,  
13'd186,  13'd264,  -13'd335,  13'd519,  13'd245,  -13'd82,  13'd671,  13'd1059,  13'd137,  13'd531,  -13'd625,  13'd1,  13'd108,  -13'd301,  13'd397,  13'd201,  
-13'd176,  13'd291,  13'd356,  -13'd534,  13'd339,  -13'd459,  13'd97,  13'd388,  -13'd235,  13'd199,  13'd194,  -13'd104,  13'd787,  -13'd566,  -13'd120,  -13'd856,  
13'd323,  13'd561,  -13'd289,  -13'd409,  13'd362,  -13'd317,  -13'd788,  13'd470,  13'd131,  13'd232,  -13'd186,  13'd518,  13'd145,  13'd256,  -13'd992,  13'd313,  
13'd725,  -13'd38,  13'd324,  13'd201,  13'd879,  13'd350,  -13'd437,  -13'd147,  -13'd344,  -13'd428,  13'd532,  -13'd94,  13'd660,  -13'd341,  13'd391,  -13'd93,  
13'd233,  13'd924,  -13'd786,  13'd532,  -13'd1121,  -13'd602,  13'd619,  13'd973,  -13'd58,  13'd47,  -13'd555,  13'd96,  13'd835,  -13'd183,  13'd183,  13'd162,  
-13'd43,  13'd236,  -13'd818,  -13'd536,  -13'd723,  -13'd292,  -13'd159,  -13'd940,  13'd478,  13'd585,  13'd134,  13'd43,  13'd103,  13'd200,  -13'd592,  13'd296,  
13'd527,  13'd83,  -13'd728,  -13'd148,  -13'd159,  -13'd199,  13'd281,  13'd609,  
-13'd284,  13'd339,  -13'd442,  13'd362,  13'd341,  13'd485,  -13'd209,  -13'd704,  13'd389,  13'd493,  13'd254,  13'd363,  13'd629,  13'd443,  -13'd503,  13'd140,  
-13'd65,  13'd381,  13'd362,  13'd758,  -13'd66,  13'd539,  -13'd390,  -13'd836,  -13'd576,  13'd723,  -13'd765,  13'd300,  -13'd192,  -13'd484,  -13'd110,  -13'd495,  
13'd213,  13'd683,  -13'd522,  13'd68,  13'd788,  13'd448,  -13'd716,  -13'd245,  -13'd491,  13'd722,  -13'd556,  13'd289,  -13'd222,  13'd400,  13'd147,  13'd51,  
13'd292,  -13'd380,  -13'd108,  13'd567,  13'd22,  13'd644,  -13'd16,  -13'd245,  -13'd55,  -13'd445,  -13'd747,  -13'd166,  13'd277,  13'd205,  13'd1055,  -13'd211,  
-13'd262,  -13'd577,  13'd114,  -13'd83,  13'd116,  13'd497,  13'd153,  13'd861,  13'd63,  -13'd370,  -13'd685,  -13'd908,  -13'd527,  -13'd403,  13'd265,  13'd993,  
13'd60,  13'd429,  13'd14,  -13'd399,  13'd185,  13'd704,  -13'd865,  13'd628,  13'd48,  -13'd757,  13'd745,  -13'd669,  13'd552,  -13'd332,  13'd337,  -13'd66,  
-13'd542,  -13'd197,  -13'd245,  13'd336,  -13'd244,  13'd790,  13'd488,  13'd746,  -13'd211,  13'd139,  -13'd509,  13'd185,  13'd174,  -13'd955,  13'd389,  13'd669,  
-13'd813,  13'd730,  13'd377,  13'd354,  -13'd27,  -13'd231,  13'd274,  13'd153,  
-13'd49,  13'd70,  -13'd1044,  13'd710,  -13'd198,  -13'd655,  13'd685,  -13'd114,  13'd91,  -13'd56,  13'd533,  13'd261,  13'd160,  13'd47,  -13'd198,  13'd512,  
-13'd226,  13'd311,  13'd458,  13'd395,  -13'd199,  13'd379,  -13'd16,  13'd150,  13'd751,  -13'd58,  13'd845,  13'd376,  13'd89,  13'd314,  13'd280,  -13'd211,  
13'd484,  -13'd0,  -13'd492,  13'd587,  -13'd567,  13'd961,  13'd421,  -13'd611,  13'd457,  13'd152,  13'd192,  13'd349,  -13'd239,  13'd159,  13'd331,  13'd856,  
-13'd147,  -13'd246,  13'd348,  -13'd385,  13'd821,  -13'd56,  13'd960,  13'd357,  13'd312,  13'd676,  -13'd669,  -13'd444,  -13'd253,  13'd799,  13'd120,  -13'd495,  
-13'd186,  -13'd251,  -13'd247,  13'd560,  13'd316,  -13'd52,  13'd121,  13'd233,  13'd308,  13'd952,  -13'd263,  -13'd427,  -13'd11,  13'd104,  -13'd305,  13'd392,  
13'd587,  13'd239,  -13'd569,  13'd794,  13'd209,  -13'd593,  13'd91,  13'd930,  13'd724,  -13'd194,  -13'd98,  13'd411,  -13'd352,  -13'd278,  -13'd162,  -13'd210,  
13'd612,  -13'd64,  -13'd398,  -13'd110,  -13'd216,  13'd15,  -13'd496,  13'd1021,  -13'd385,  13'd535,  13'd257,  13'd283,  13'd440,  -13'd324,  13'd729,  -13'd182,  
-13'd367,  13'd103,  -13'd93,  13'd353,  13'd683,  -13'd146,  13'd436,  -13'd190,  
-13'd1204,  13'd253,  13'd439,  -13'd85,  -13'd1114,  13'd521,  13'd100,  -13'd272,  -13'd792,  -13'd779,  13'd575,  -13'd353,  -13'd600,  13'd38,  13'd329,  13'd253,  
-13'd730,  13'd127,  13'd177,  13'd170,  13'd337,  -13'd167,  13'd162,  -13'd644,  -13'd325,  13'd38,  13'd645,  13'd538,  -13'd87,  13'd500,  -13'd72,  -13'd426,  
-13'd462,  13'd68,  -13'd530,  13'd33,  13'd1272,  13'd475,  -13'd905,  13'd93,  13'd115,  13'd237,  13'd98,  -13'd40,  -13'd346,  13'd179,  13'd87,  13'd11,  
13'd207,  -13'd533,  13'd751,  -13'd636,  13'd270,  13'd15,  -13'd239,  13'd52,  -13'd1254,  13'd442,  13'd815,  -13'd286,  -13'd353,  -13'd242,  13'd897,  13'd316,  
13'd639,  13'd117,  13'd618,  -13'd372,  -13'd61,  -13'd6,  13'd184,  13'd109,  13'd455,  -13'd1209,  13'd285,  13'd362,  -13'd14,  -13'd439,  -13'd163,  -13'd93,  
13'd33,  13'd488,  -13'd315,  -13'd650,  13'd705,  13'd693,  13'd609,  13'd308,  13'd403,  13'd22,  13'd458,  -13'd405,  -13'd4,  -13'd91,  13'd99,  13'd806,  
13'd456,  13'd82,  13'd319,  -13'd791,  13'd340,  -13'd772,  13'd600,  13'd196,  13'd137,  -13'd416,  -13'd210,  -13'd505,  -13'd123,  13'd1849,  -13'd639,  13'd224,  
-13'd468,  -13'd204,  -13'd103,  13'd48,  13'd110,  -13'd54,  -13'd524,  13'd794,  
-13'd1241,  13'd220,  -13'd273,  -13'd35,  13'd60,  13'd221,  13'd711,  13'd27,  13'd1118,  13'd31,  13'd916,  13'd161,  13'd749,  13'd186,  -13'd308,  13'd64,  
-13'd551,  -13'd11,  13'd674,  13'd759,  -13'd396,  13'd815,  -13'd524,  -13'd674,  -13'd307,  -13'd187,  13'd100,  13'd610,  -13'd126,  13'd50,  13'd355,  -13'd660,  
-13'd443,  -13'd237,  -13'd203,  13'd630,  -13'd346,  -13'd53,  13'd340,  -13'd69,  -13'd168,  13'd507,  -13'd693,  -13'd15,  -13'd429,  13'd109,  13'd389,  13'd1077,  
-13'd285,  13'd178,  13'd696,  -13'd194,  -13'd365,  -13'd481,  -13'd207,  -13'd235,  -13'd337,  13'd170,  13'd94,  -13'd585,  13'd469,  -13'd108,  13'd628,  13'd111,  
-13'd393,  13'd71,  13'd184,  13'd865,  13'd96,  13'd466,  13'd350,  13'd439,  13'd234,  -13'd530,  13'd48,  13'd119,  -13'd729,  13'd348,  -13'd529,  13'd365,  
13'd419,  13'd236,  -13'd56,  13'd87,  13'd365,  13'd198,  13'd598,  13'd178,  -13'd117,  13'd361,  13'd31,  13'd465,  -13'd141,  13'd128,  -13'd5,  -13'd176,  
13'd129,  13'd450,  -13'd94,  13'd80,  -13'd788,  13'd219,  -13'd316,  13'd828,  -13'd382,  13'd654,  -13'd66,  -13'd373,  -13'd575,  13'd1085,  -13'd169,  13'd82,  
-13'd121,  -13'd507,  13'd890,  13'd663,  -13'd376,  13'd218,  -13'd323,  -13'd57,  
13'd467,  -13'd176,  13'd499,  13'd297,  13'd263,  -13'd437,  -13'd342,  -13'd307,  -13'd69,  13'd295,  -13'd105,  -13'd846,  13'd703,  13'd361,  13'd657,  13'd0,  
-13'd89,  13'd184,  -13'd50,  -13'd288,  13'd504,  -13'd21,  -13'd513,  13'd266,  13'd226,  13'd45,  -13'd197,  -13'd478,  13'd533,  13'd447,  13'd632,  13'd813,  
13'd70,  13'd113,  -13'd505,  -13'd119,  13'd630,  13'd220,  13'd905,  -13'd924,  -13'd361,  13'd648,  -13'd208,  -13'd197,  -13'd276,  13'd60,  -13'd741,  -13'd522,  
-13'd149,  13'd412,  13'd93,  13'd18,  13'd805,  13'd502,  -13'd770,  13'd378,  13'd203,  -13'd658,  13'd166,  13'd260,  13'd304,  13'd81,  -13'd422,  -13'd498,  
13'd738,  13'd79,  13'd129,  -13'd170,  -13'd306,  13'd587,  13'd469,  -13'd124,  13'd52,  -13'd401,  13'd267,  -13'd519,  13'd76,  13'd518,  -13'd372,  -13'd13,  
13'd160,  -13'd158,  -13'd487,  13'd1142,  13'd581,  -13'd16,  13'd164,  13'd173,  -13'd820,  -13'd200,  -13'd13,  -13'd883,  13'd252,  13'd401,  -13'd380,  -13'd648,  
-13'd202,  13'd250,  -13'd570,  -13'd42,  -13'd570,  13'd406,  -13'd129,  13'd311,  -13'd666,  13'd618,  -13'd62,  13'd718,  -13'd358,  -13'd151,  13'd684,  13'd283,  
-13'd69,  -13'd109,  13'd187,  -13'd18,  -13'd14,  13'd134,  -13'd118,  -13'd20,  
-13'd947,  -13'd685,  13'd929,  -13'd357,  -13'd425,  -13'd405,  -13'd71,  13'd815,  13'd21,  13'd427,  13'd1382,  13'd9,  -13'd286,  13'd468,  -13'd656,  13'd605,  
-13'd693,  13'd289,  13'd591,  -13'd552,  -13'd242,  -13'd99,  -13'd4,  13'd122,  13'd565,  13'd355,  13'd295,  13'd326,  -13'd336,  -13'd172,  -13'd619,  13'd171,  
13'd448,  13'd455,  -13'd194,  13'd363,  13'd89,  13'd738,  -13'd337,  13'd753,  -13'd64,  13'd681,  13'd384,  13'd563,  13'd685,  13'd552,  -13'd131,  13'd100,  
-13'd260,  13'd414,  13'd531,  13'd317,  13'd85,  -13'd869,  13'd214,  13'd688,  13'd408,  -13'd588,  13'd586,  13'd461,  -13'd374,  -13'd168,  13'd374,  13'd831,  
13'd110,  13'd376,  -13'd0,  -13'd59,  -13'd289,  -13'd251,  13'd347,  -13'd95,  -13'd2,  -13'd124,  13'd140,  -13'd308,  -13'd164,  -13'd544,  13'd460,  -13'd173,  
-13'd430,  -13'd204,  13'd76,  -13'd469,  13'd362,  13'd17,  -13'd61,  13'd137,  13'd629,  13'd185,  13'd556,  13'd285,  -13'd634,  13'd75,  -13'd189,  13'd412,  
13'd10,  13'd863,  13'd246,  13'd301,  -13'd146,  -13'd64,  -13'd329,  13'd726,  13'd433,  -13'd299,  -13'd416,  -13'd340,  13'd373,  13'd915,  -13'd87,  -13'd284,  
13'd347,  -13'd516,  -13'd309,  13'd94,  13'd221,  -13'd88,  -13'd165,  13'd557,  
13'd379,  -13'd427,  -13'd179,  13'd45,  13'd266,  -13'd468,  -13'd400,  13'd418,  -13'd227,  13'd299,  -13'd1019,  13'd228,  13'd98,  -13'd14,  13'd643,  -13'd743,  
13'd128,  -13'd107,  -13'd1389,  -13'd214,  13'd561,  -13'd170,  -13'd308,  -13'd516,  -13'd566,  13'd243,  13'd66,  -13'd656,  -13'd228,  13'd807,  13'd314,  -13'd88,  
13'd467,  13'd713,  -13'd304,  13'd477,  13'd479,  13'd256,  -13'd526,  -13'd927,  13'd79,  13'd161,  13'd356,  -13'd1403,  13'd732,  13'd55,  -13'd565,  -13'd577,  
-13'd552,  -13'd238,  13'd713,  -13'd939,  -13'd501,  13'd787,  -13'd209,  13'd330,  -13'd538,  -13'd32,  -13'd893,  13'd431,  -13'd388,  -13'd709,  13'd436,  13'd120,  
13'd76,  13'd277,  -13'd145,  -13'd459,  -13'd618,  13'd34,  13'd385,  -13'd397,  -13'd400,  13'd288,  13'd162,  13'd208,  13'd72,  13'd506,  13'd205,  13'd211,  
13'd266,  -13'd877,  -13'd487,  -13'd138,  13'd362,  13'd30,  13'd75,  13'd291,  -13'd993,  13'd201,  13'd240,  -13'd843,  -13'd49,  13'd666,  -13'd646,  13'd356,  
-13'd220,  13'd322,  -13'd145,  -13'd649,  13'd764,  -13'd89,  -13'd188,  13'd315,  -13'd96,  -13'd202,  -13'd505,  -13'd248,  -13'd431,  13'd10,  -13'd165,  13'd887,  
-13'd652,  13'd501,  13'd155,  13'd265,  -13'd500,  -13'd452,  13'd301,  -13'd100,  
13'd117,  -13'd409,  13'd523,  -13'd17,  13'd169,  13'd60,  13'd359,  -13'd115,  13'd213,  -13'd440,  13'd120,  13'd205,  -13'd722,  13'd111,  -13'd552,  -13'd539,  
13'd567,  13'd438,  13'd593,  13'd419,  -13'd392,  -13'd60,  13'd250,  -13'd83,  13'd633,  13'd282,  -13'd395,  -13'd250,  -13'd66,  13'd600,  -13'd627,  -13'd817,  
-13'd78,  13'd77,  13'd154,  13'd69,  -13'd472,  13'd562,  13'd69,  13'd699,  13'd266,  13'd150,  13'd460,  -13'd436,  -13'd414,  -13'd20,  13'd111,  13'd704,  
13'd8,  13'd322,  -13'd462,  13'd389,  -13'd1005,  -13'd281,  13'd840,  -13'd533,  13'd236,  13'd413,  13'd25,  -13'd460,  13'd162,  -13'd561,  -13'd16,  -13'd355,  
-13'd267,  13'd299,  13'd62,  -13'd275,  13'd314,  13'd396,  13'd72,  13'd252,  -13'd146,  13'd37,  13'd5,  -13'd826,  13'd59,  13'd282,  -13'd65,  -13'd697,  
-13'd272,  -13'd535,  13'd628,  13'd884,  13'd585,  13'd383,  -13'd189,  -13'd586,  13'd603,  13'd626,  13'd477,  -13'd143,  -13'd762,  13'd906,  -13'd367,  13'd603,  
-13'd288,  -13'd223,  13'd537,  13'd499,  -13'd55,  13'd54,  13'd341,  13'd903,  -13'd233,  13'd39,  -13'd194,  13'd313,  13'd217,  -13'd841,  13'd867,  -13'd633,  
-13'd705,  -13'd513,  13'd102,  13'd139,  13'd366,  -13'd182,  -13'd149,  -13'd274,  
-13'd329,  13'd447,  -13'd955,  13'd552,  13'd221,  -13'd76,  -13'd62,  13'd81,  13'd115,  -13'd541,  -13'd867,  13'd483,  13'd893,  -13'd510,  -13'd346,  13'd2,  
-13'd88,  13'd32,  -13'd83,  -13'd42,  -13'd85,  13'd58,  13'd45,  -13'd110,  -13'd174,  -13'd830,  13'd415,  13'd115,  13'd119,  -13'd304,  13'd664,  -13'd755,  
-13'd213,  -13'd364,  -13'd188,  13'd330,  -13'd748,  13'd179,  13'd693,  -13'd147,  13'd421,  -13'd286,  -13'd659,  13'd148,  13'd238,  -13'd423,  13'd264,  13'd773,  
-13'd490,  -13'd1146,  -13'd144,  -13'd333,  13'd514,  13'd545,  -13'd795,  -13'd91,  13'd573,  13'd231,  -13'd244,  -13'd779,  13'd1010,  -13'd154,  13'd193,  -13'd168,  
13'd25,  13'd65,  -13'd384,  -13'd167,  13'd739,  -13'd233,  13'd247,  13'd779,  -13'd388,  13'd495,  -13'd152,  13'd779,  13'd391,  13'd722,  -13'd596,  -13'd182,  
13'd408,  13'd629,  -13'd768,  13'd364,  -13'd619,  13'd29,  13'd384,  13'd706,  13'd176,  13'd34,  13'd47,  13'd188,  -13'd185,  -13'd0,  -13'd361,  13'd832,  
-13'd172,  13'd72,  13'd466,  13'd663,  13'd87,  -13'd284,  13'd604,  13'd807,  -13'd315,  -13'd128,  13'd228,  13'd985,  13'd152,  -13'd34,  13'd442,  13'd283,  
-13'd76,  13'd881,  13'd515,  13'd104,  13'd769,  -13'd638,  13'd97,  -13'd148
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule


module bias_fc3_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC3-1][0:`OUTPUT_NUM_FC3-1][`WD_BIAS:0] weight	 = {
-24'd186531,  24'd166143,  -24'd211411,  -24'd80228,  -24'd155665,  24'd207658,  -24'd315652,  -24'd209780,  24'd326774,  24'd153726
	};

	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule




module wieght_fc3_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3*`OUTPUT_BATCH_FC3)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC2*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC3*`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3-1][0:`OUTPUT_NUM_FC3-1][0:`OUTPUT_NUM_FC2-1][`WD:0] weight	 = {
-13'd49,  13'd427,  -13'd64,  -13'd126,  13'd141,  13'd229,  13'd119,  -13'd109,  -13'd464,  -13'd361,  13'd1021,  -13'd690,  -13'd227,  -13'd39,  -13'd512,  13'd408,  
13'd592,  13'd95,  -13'd96,  13'd1043,  13'd1297,  -13'd979,  -13'd686,  -13'd88,  -13'd807,  13'd655,  13'd250,  -13'd77,  -13'd372,  13'd499,  13'd170,  13'd617,  
-13'd587,  -13'd989,  -13'd343,  -13'd942,  -13'd263,  13'd351,  13'd252,  -13'd258,  13'd386,  -13'd71,  13'd730,  -13'd341,  -13'd877,  13'd176,  -13'd183,  13'd164,  
-13'd1023,  -13'd133,  13'd597,  13'd161,  13'd1023,  -13'd362,  -13'd630,  13'd578,  -13'd376,  13'd1034,  13'd2,  -13'd130,  -13'd234,  -13'd241,  13'd183,  -13'd579,  
13'd857,  -13'd914,  -13'd242,  -13'd175,  -13'd464,  -13'd511,  -13'd38,  -13'd1220,  -13'd56,  -13'd273,  -13'd465,  13'd150,  13'd97,  -13'd356,  13'd601,  -13'd196,  
-13'd236,  -13'd585,  13'd776,  -13'd523,  
13'd570,  -13'd855,  13'd166,  -13'd396,  -13'd57,  13'd211,  13'd429,  -13'd324,  -13'd73,  -13'd522,  -13'd961,  13'd479,  13'd59,  13'd689,  13'd253,  13'd249,  
-13'd579,  13'd525,  -13'd517,  -13'd397,  13'd890,  -13'd274,  -13'd26,  13'd71,  -13'd875,  -13'd100,  -13'd169,  13'd658,  13'd497,  -13'd102,  13'd675,  -13'd227,  
13'd9,  -13'd536,  -13'd4,  13'd804,  -13'd450,  -13'd493,  -13'd255,  -13'd788,  13'd608,  -13'd387,  -13'd1149,  -13'd868,  13'd560,  13'd392,  -13'd3,  13'd392,  
-13'd427,  13'd693,  -13'd979,  -13'd432,  -13'd136,  13'd401,  13'd1044,  -13'd494,  -13'd261,  -13'd316,  -13'd1157,  13'd1007,  -13'd510,  13'd120,  -13'd712,  -13'd226,  
13'd786,  -13'd472,  13'd256,  13'd1119,  13'd368,  -13'd733,  -13'd501,  13'd622,  13'd465,  13'd130,  -13'd803,  -13'd450,  -13'd47,  -13'd844,  -13'd702,  13'd256,  
13'd425,  -13'd1007,  13'd1005,  -13'd157,  
-13'd707,  -13'd718,  13'd458,  -13'd97,  13'd966,  13'd395,  -13'd396,  13'd95,  13'd270,  -13'd384,  13'd467,  13'd848,  13'd157,  -13'd666,  -13'd244,  -13'd318,  
-13'd138,  -13'd1261,  -13'd659,  13'd418,  13'd798,  13'd108,  -13'd324,  -13'd677,  13'd53,  -13'd214,  -13'd87,  -13'd246,  -13'd386,  13'd746,  -13'd1326,  -13'd55,  
-13'd1235,  -13'd243,  13'd53,  -13'd659,  13'd170,  13'd576,  13'd196,  13'd905,  -13'd54,  -13'd189,  13'd188,  -13'd408,  13'd56,  -13'd101,  13'd462,  13'd411,  
13'd525,  13'd598,  -13'd1123,  -13'd868,  -13'd257,  -13'd297,  -13'd424,  -13'd342,  13'd167,  13'd603,  13'd15,  13'd213,  -13'd71,  -13'd843,  -13'd63,  13'd640,  
13'd293,  -13'd653,  13'd209,  -13'd485,  -13'd280,  13'd316,  13'd299,  13'd177,  -13'd573,  13'd352,  -13'd470,  13'd82,  -13'd188,  13'd850,  13'd216,  -13'd644,  
13'd946,  -13'd202,  -13'd53,  -13'd486,  
-13'd5,  -13'd446,  13'd66,  -13'd958,  13'd553,  13'd84,  -13'd493,  -13'd423,  13'd172,  -13'd300,  -13'd642,  -13'd500,  13'd951,  -13'd572,  -13'd567,  13'd179,  
-13'd558,  13'd283,  -13'd382,  13'd757,  -13'd1263,  -13'd506,  -13'd557,  -13'd750,  -13'd59,  13'd204,  -13'd603,  13'd188,  -13'd661,  13'd480,  -13'd130,  -13'd188,  
13'd68,  13'd255,  -13'd544,  13'd505,  13'd291,  -13'd449,  -13'd174,  13'd496,  -13'd431,  -13'd220,  13'd666,  13'd323,  13'd564,  -13'd788,  -13'd296,  -13'd485,  
13'd604,  -13'd945,  13'd101,  13'd697,  -13'd661,  -13'd19,  -13'd235,  -13'd383,  -13'd404,  -13'd348,  13'd458,  13'd33,  13'd88,  13'd143,  -13'd76,  13'd228,  
-13'd766,  13'd1297,  -13'd130,  13'd343,  13'd22,  13'd21,  -13'd793,  13'd614,  -13'd930,  13'd410,  -13'd284,  13'd9,  13'd576,  13'd62,  13'd4,  -13'd238,  
-13'd886,  -13'd233,  13'd141,  13'd1023,  
-13'd592,  13'd656,  13'd31,  13'd226,  -13'd644,  13'd387,  13'd1039,  13'd555,  -13'd812,  -13'd8,  -13'd290,  -13'd493,  -13'd331,  13'd735,  13'd416,  -13'd747,  
13'd716,  -13'd413,  -13'd976,  -13'd149,  -13'd663,  13'd348,  -13'd100,  -13'd1016,  13'd423,  -13'd206,  -13'd1518,  -13'd236,  13'd844,  13'd312,  -13'd789,  -13'd633,  
13'd15,  -13'd836,  -13'd200,  13'd73,  -13'd670,  13'd442,  13'd534,  -13'd886,  13'd5,  -13'd256,  13'd53,  13'd854,  13'd208,  13'd511,  -13'd148,  13'd186,  
13'd398,  -13'd266,  13'd443,  -13'd420,  13'd491,  13'd4,  -13'd352,  -13'd172,  -13'd121,  13'd191,  -13'd354,  13'd802,  -13'd38,  -13'd145,  -13'd622,  13'd588,  
13'd209,  -13'd803,  13'd78,  13'd794,  -13'd981,  -13'd482,  13'd679,  -13'd452,  -13'd890,  -13'd713,  13'd480,  13'd700,  -13'd821,  13'd462,  -13'd847,  13'd642,  
-13'd641,  13'd464,  -13'd539,  -13'd635,  
13'd1113,  13'd558,  -13'd739,  -13'd738,  13'd1013,  -13'd627,  -13'd768,  13'd252,  13'd588,  13'd603,  13'd230,  13'd1022,  -13'd695,  -13'd593,  13'd89,  -13'd360,  
13'd295,  13'd752,  13'd426,  13'd413,  -13'd615,  13'd320,  -13'd462,  13'd673,  13'd627,  13'd348,  13'd450,  13'd100,  -13'd342,  13'd28,  13'd225,  -13'd320,  
-13'd13,  -13'd118,  13'd285,  13'd1075,  -13'd610,  -13'd1128,  -13'd910,  13'd259,  13'd408,  13'd32,  -13'd677,  -13'd561,  -13'd665,  -13'd446,  -13'd316,  13'd0,  
13'd618,  13'd677,  13'd87,  13'd616,  13'd238,  -13'd905,  -13'd1028,  13'd257,  -13'd345,  -13'd217,  13'd272,  -13'd699,  13'd3,  13'd27,  13'd46,  -13'd767,  
-13'd45,  -13'd180,  13'd682,  13'd178,  -13'd87,  -13'd450,  -13'd332,  -13'd71,  13'd1019,  -13'd84,  13'd568,  13'd259,  13'd254,  -13'd193,  13'd24,  13'd542,  
-13'd750,  13'd337,  -13'd718,  13'd162,  
13'd927,  -13'd505,  -13'd112,  -13'd29,  -13'd47,  -13'd652,  -13'd114,  13'd548,  13'd206,  13'd556,  -13'd392,  -13'd562,  -13'd1515,  -13'd87,  -13'd610,  -13'd587,  
13'd571,  -13'd218,  -13'd761,  -13'd520,  13'd167,  13'd176,  -13'd724,  -13'd357,  13'd377,  -13'd306,  -13'd28,  13'd21,  -13'd848,  13'd99,  13'd555,  13'd355,  
-13'd346,  13'd870,  -13'd63,  -13'd261,  -13'd742,  -13'd640,  13'd403,  -13'd409,  -13'd318,  -13'd735,  13'd1085,  -13'd905,  13'd75,  -13'd279,  13'd393,  -13'd60,  
-13'd259,  -13'd783,  13'd532,  -13'd479,  13'd49,  13'd452,  13'd134,  13'd385,  -13'd1,  13'd200,  13'd313,  -13'd12,  13'd323,  -13'd717,  13'd328,  -13'd932,  
13'd278,  13'd462,  -13'd129,  13'd50,  -13'd53,  13'd207,  13'd319,  -13'd516,  13'd489,  -13'd352,  13'd222,  -13'd711,  -13'd540,  13'd324,  -13'd500,  13'd125,  
13'd264,  13'd403,  -13'd406,  -13'd1225,  
-13'd706,  -13'd163,  13'd344,  -13'd1349,  -13'd551,  13'd350,  -13'd1131,  -13'd344,  -13'd439,  -13'd379,  -13'd1128,  13'd224,  13'd169,  13'd314,  -13'd478,  13'd66,  
13'd450,  -13'd45,  -13'd464,  -13'd302,  -13'd266,  -13'd340,  -13'd426,  -13'd398,  -13'd214,  -13'd89,  -13'd107,  -13'd378,  13'd907,  -13'd197,  13'd303,  -13'd45,  
13'd21,  -13'd177,  13'd1116,  -13'd356,  13'd128,  13'd838,  -13'd676,  -13'd251,  -13'd279,  13'd165,  -13'd1130,  -13'd31,  13'd815,  13'd830,  -13'd339,  -13'd157,  
13'd122,  13'd220,  13'd333,  -13'd770,  13'd380,  13'd133,  13'd74,  -13'd564,  13'd313,  -13'd1313,  -13'd765,  13'd481,  -13'd98,  13'd672,  -13'd505,  -13'd490,  
-13'd117,  13'd1044,  13'd31,  -13'd1187,  13'd732,  -13'd324,  13'd93,  13'd36,  13'd117,  -13'd117,  13'd325,  13'd136,  13'd517,  13'd412,  13'd534,  -13'd41,  
13'd349,  -13'd762,  13'd174,  13'd4,  
13'd51,  13'd524,  13'd387,  -13'd111,  -13'd18,  -13'd29,  13'd6,  -13'd417,  -13'd136,  13'd1044,  -13'd847,  -13'd1005,  13'd121,  -13'd786,  -13'd41,  13'd134,  
13'd235,  13'd308,  13'd489,  13'd129,  13'd69,  13'd591,  -13'd99,  -13'd380,  13'd60,  -13'd465,  -13'd751,  13'd84,  -13'd568,  -13'd400,  -13'd1110,  -13'd481,  
-13'd734,  13'd463,  -13'd404,  13'd446,  13'd129,  13'd75,  -13'd122,  13'd286,  -13'd76,  13'd123,  -13'd509,  13'd941,  -13'd704,  13'd650,  13'd125,  13'd143,  
-13'd672,  -13'd946,  -13'd638,  13'd580,  13'd529,  13'd520,  13'd322,  13'd260,  -13'd144,  -13'd606,  13'd169,  -13'd634,  13'd695,  -13'd629,  13'd569,  -13'd1,  
13'd477,  13'd604,  -13'd621,  -13'd384,  13'd26,  -13'd884,  -13'd781,  13'd8,  13'd421,  13'd47,  13'd271,  -13'd926,  -13'd626,  13'd79,  13'd169,  -13'd959,  
13'd632,  13'd898,  -13'd29,  -13'd175,  
13'd196,  13'd252,  13'd373,  13'd200,  13'd355,  -13'd432,  13'd337,  13'd295,  -13'd393,  -13'd551,  13'd325,  13'd415,  13'd623,  13'd695,  13'd404,  13'd213,  
-13'd802,  -13'd66,  -13'd225,  -13'd354,  -13'd10,  -13'd379,  13'd538,  13'd133,  13'd591,  -13'd202,  13'd218,  -13'd293,  13'd294,  -13'd1145,  -13'd561,  -13'd240,  
13'd103,  -13'd728,  13'd202,  -13'd88,  -13'd410,  13'd817,  13'd302,  13'd632,  13'd707,  13'd638,  -13'd287,  13'd135,  13'd369,  -13'd124,  13'd148,  -13'd69,  
-13'd1144,  -13'd366,  -13'd96,  13'd408,  13'd442,  -13'd82,  -13'd1321,  -13'd66,  -13'd132,  13'd555,  13'd340,  -13'd971,  13'd95,  13'd473,  13'd1148,  13'd570,  
-13'd241,  -13'd1477,  13'd271,  13'd123,  -13'd12,  13'd775,  13'd658,  13'd510,  -13'd284,  -13'd1319,  13'd650,  -13'd838,  -13'd121,  -13'd924,  -13'd664,  13'd221,  
-13'd814,  -13'd664,  -13'd285,  -13'd22
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule

