// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION
`include "global.v"


module bias_conv1_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV1-1][0:`OUTPUT_NUM_CONV1-1][`WD_BIAS:0] weight	 = {	
		-24'd33091,  -24'd345382,  -24'd986031,  -24'd314271,  24'd400309,  -24'd448129
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_conv1_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV1*`KERNEL_SIZE_CONV1-1][0:`OUTPUT_NUM_CONV1-1][11:0] weight	 = {
12'd61,  12'd116,  -12'd227,  12'd222,  -12'd397,  -12'd767,  
12'd237,  -12'd190,  -12'd129,  -12'd85,  -12'd493,  -12'd470,  
-12'd486,  -12'd341,  -12'd92,  12'd128,  -12'd690,  12'd17,  
-12'd479,  -12'd93,  12'd228,  12'd266,  -12'd537,  12'd214,  
-12'd784,  12'd252,  12'd61,  -12'd166,  -12'd564,  12'd590,  

12'd422,  -12'd194,  -12'd322,  12'd524,  -12'd44,  -12'd551,  
12'd52,  -12'd288,  -12'd104,  12'd256,  -12'd735,  12'd177,  
12'd231,  12'd25,  12'd254,  12'd349,  -12'd443,  12'd325,  
-12'd310,  12'd240,  12'd395,  12'd476,  -12'd249,  12'd531,  
-12'd697,  12'd0,  12'd155,  -12'd332,  -12'd452,  -12'd167,  

12'd221,  -12'd96,  -12'd423,  12'd429,  12'd88,  -12'd208,  
12'd637,  12'd53,  12'd246,  12'd222,  12'd186,  12'd177,  
12'd640,  -12'd64,  12'd357,  12'd338,  12'd104,  12'd512,  
12'd194,  12'd438,  12'd489,  12'd374,  12'd124,  12'd244,  
12'd313,  12'd279,  -12'd145,  12'd79,  12'd478,  -12'd518,  

-12'd433,  -12'd94,  -12'd51,  -12'd1,  12'd661,  12'd40,  
12'd367,  12'd87,  12'd131,  12'd326,  12'd635,  12'd259,  
12'd18,  12'd560,  12'd745,  12'd419,  12'd483,  12'd442,  
12'd531,  12'd505,  12'd42,  12'd602,  12'd575,  -12'd27,  
12'd180,  -12'd147,  -12'd350,  12'd577,  12'd311,  -12'd895,  

-12'd381,  12'd20,  12'd465,  12'd1,  12'd426,  12'd110,  
-12'd265,  12'd277,  12'd361,  -12'd445,  12'd116,  12'd8,  
-12'd183,  12'd13,  12'd333,  -12'd4,  12'd344,  12'd306,  
12'd287,  12'd512,  -12'd208,  12'd100,  -12'd55,  -12'd54,  
-12'd110,  12'd365,  -12'd314,  12'd492,  12'd108,  -12'd470
		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule	


module bias_conv2_rom(
	input							clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_CONV2-1][0:`OUTPUT_NUM_CONV2-1][`WD_BIAS:0] weight	 = {
	-24'd492928,  -24'd252352,  24'd425549,  -24'd126681,  -24'd362367,  -24'd84127,  24'd122339,  -24'd193094,  24'd178645,  24'd56283,  -24'd15047,  -24'd647019,  -24'd375850,  24'd168062,  -24'd242871,  -24'd1026233		};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule



module wieght_conv2_rom(
	input			clk,
	input			rstn,
	input	[9:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV1*`OUTPUT_NUM_CONV2 -1:0]	qa
	);
	
	
	logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][`WD:0] weight	 = {
12'd233,  -12'd130,  12'd265,  12'd126,  -12'd78,  12'd263,  
-12'd355,  -12'd267,  12'd203,  12'd114,  -12'd221,  -12'd269,  
12'd319,  -12'd352,  -12'd489,  -12'd262,  -12'd3,  12'd107,  
-12'd14,  12'd100,  -12'd369,  -12'd124,  -12'd204,  -12'd557,  
12'd118,  -12'd340,  -12'd113,  -12'd348,  -12'd311,  12'd61,  
-12'd363,  -12'd207,  12'd140,  -12'd55,  -12'd198,  12'd214,  
12'd68,  12'd87,  -12'd205,  12'd250,  -12'd159,  12'd63,  
12'd31,  12'd14,  -12'd310,  12'd67,  -12'd348,  12'd74,  
12'd61,  -12'd541,  -12'd311,  -12'd153,  12'd193,  -12'd246,  
12'd370,  -12'd493,  -12'd491,  -12'd6,  -12'd713,  12'd274,  
-12'd267,  -12'd160,  -12'd19,  -12'd75,  -12'd30,  -12'd546,  
-12'd179,  -12'd146,  -12'd322,  -12'd1,  12'd114,  12'd92,  
-12'd108,  -12'd223,  -12'd109,  -12'd123,  12'd56,  12'd206,  
12'd300,  12'd65,  -12'd157,  12'd464,  12'd31,  -12'd70,  
12'd30,  12'd229,  -12'd144,  12'd141,  12'd300,  -12'd333,  
-12'd171,  12'd121,  -12'd78,  -12'd74,  -12'd178,  -12'd9,  

-12'd140,  12'd11,  -12'd253,  -12'd381,  -12'd114,  -12'd159,  
12'd136,  -12'd140,  -12'd154,  12'd353,  -12'd214,  -12'd232,  
-12'd671,  -12'd369,  -12'd12,  -12'd379,  -12'd192,  -12'd127,  
12'd85,  12'd28,  -12'd147,  -12'd281,  -12'd31,  12'd133,  
-12'd516,  -12'd62,  12'd222,  -12'd91,  -12'd286,  12'd207,  
-12'd81,  12'd271,  -12'd133,  12'd36,  -12'd73,  -12'd362,  
-12'd290,  12'd274,  -12'd115,  12'd353,  -12'd51,  12'd297,  
-12'd142,  -12'd147,  -12'd258,  12'd171,  -12'd12,  12'd60,  
-12'd136,  -12'd97,  12'd76,  -12'd272,  12'd16,  -12'd259,  
-12'd20,  -12'd506,  12'd302,  -12'd14,  -12'd495,  12'd77,  
-12'd112,  -12'd205,  12'd135,  -12'd135,  12'd438,  12'd29,  
-12'd440,  -12'd5,  -12'd369,  12'd172,  12'd127,  -12'd17,  
12'd255,  -12'd46,  12'd121,  -12'd392,  -12'd56,  -12'd357,  
-12'd33,  -12'd408,  12'd316,  -12'd26,  12'd325,  -12'd28,  
12'd165,  12'd97,  12'd347,  -12'd15,  12'd116,  -12'd329,  
-12'd145,  12'd244,  -12'd76,  -12'd63,  12'd21,  -12'd231,  

-12'd8,  -12'd116,  12'd46,  -12'd372,  -12'd67,  -12'd297,  
12'd335,  -12'd299,  -12'd247,  12'd118,  -12'd80,  12'd50,  
-12'd259,  -12'd115,  -12'd302,  12'd399,  -12'd443,  -12'd300,  
12'd158,  -12'd57,  12'd141,  -12'd207,  -12'd12,  12'd355,  
-12'd134,  -12'd208,  12'd58,  12'd43,  -12'd716,  -12'd131,  
12'd307,  12'd158,  12'd27,  12'd88,  -12'd79,  -12'd449,  
12'd74,  -12'd289,  -12'd14,  -12'd275,  12'd298,  12'd122,  
-12'd190,  12'd241,  12'd302,  12'd77,  -12'd290,  12'd175,  
-12'd291,  -12'd52,  -12'd303,  -12'd196,  -12'd253,  -12'd291,  
-12'd71,  -12'd403,  -12'd237,  -12'd184,  -12'd616,  12'd203,  
12'd144,  12'd84,  -12'd173,  -12'd160,  12'd239,  -12'd460,  
12'd311,  -12'd245,  -12'd260,  12'd159,  12'd399,  -12'd219,  
-12'd314,  -12'd72,  -12'd275,  -12'd148,  -12'd5,  -12'd51,  
-12'd131,  -12'd117,  -12'd155,  -12'd150,  -12'd289,  -12'd308,  
-12'd29,  12'd288,  -12'd141,  12'd73,  12'd599,  -12'd196,  
-12'd1,  12'd85,  -12'd15,  12'd286,  12'd178,  -12'd727,  

12'd600,  -12'd248,  -12'd345,  -12'd76,  -12'd226,  -12'd494,  
12'd112,  12'd338,  -12'd198,  12'd229,  -12'd148,  -12'd172,  
12'd165,  12'd73,  12'd240,  12'd98,  -12'd489,  12'd145,  
-12'd353,  -12'd410,  -12'd153,  -12'd418,  -12'd203,  12'd321,  
12'd219,  12'd39,  -12'd247,  12'd165,  -12'd638,  -12'd515,  
12'd126,  -12'd107,  -12'd74,  -12'd222,  12'd341,  -12'd417,  
-12'd186,  -12'd50,  -12'd93,  12'd128,  12'd156,  12'd257,  
12'd31,  -12'd149,  -12'd117,  12'd13,  -12'd107,  12'd328,  
-12'd9,  -12'd5,  -12'd34,  -12'd508,  12'd253,  12'd173,  
-12'd91,  -12'd97,  12'd289,  -12'd299,  -12'd605,  -12'd97,  
-12'd114,  12'd115,  12'd299,  -12'd39,  12'd158,  12'd67,  
12'd91,  -12'd214,  -12'd265,  12'd349,  -12'd87,  -12'd628,  
-12'd269,  12'd73,  12'd156,  -12'd213,  -12'd11,  12'd16,  
-12'd489,  -12'd17,  -12'd114,  -12'd196,  -12'd541,  -12'd288,  
-12'd62,  -12'd340,  -12'd104,  -12'd221,  12'd191,  -12'd238,  
12'd145,  12'd381,  -12'd217,  -12'd120,  12'd455,  -12'd166,  

12'd337,  -12'd13,  12'd167,  -12'd14,  12'd17,  12'd266,  
12'd354,  12'd52,  12'd26,  -12'd170,  12'd473,  -12'd13,  
-12'd43,  -12'd261,  12'd108,  12'd91,  -12'd187,  12'd230,  
-12'd195,  -12'd59,  12'd89,  -12'd250,  12'd21,  12'd298,  
12'd539,  12'd168,  -12'd135,  12'd666,  12'd425,  12'd82,  
-12'd113,  -12'd239,  -12'd152,  -12'd754,  -12'd150,  12'd269,  
-12'd364,  -12'd307,  -12'd165,  12'd268,  -12'd111,  12'd573,  
12'd69,  -12'd38,  -12'd213,  12'd58,  -12'd257,  -12'd38,  
-12'd154,  12'd233,  -12'd65,  -12'd213,  12'd139,  -12'd97,  
-12'd331,  12'd266,  12'd231,  12'd340,  -12'd214,  -12'd235,  
-12'd221,  12'd102,  12'd162,  12'd110,  -12'd220,  -12'd72,  
12'd357,  -12'd294,  -12'd490,  -12'd397,  12'd146,  -12'd710,  
-12'd46,  12'd183,  12'd239,  12'd193,  -12'd224,  -12'd104,  
12'd332,  12'd309,  12'd433,  -12'd152,  -12'd456,  12'd487,  
-12'd99,  -12'd259,  12'd15,  -12'd178,  12'd348,  12'd31,  
-12'd76,  12'd94,  12'd82,  12'd19,  12'd334,  -12'd180,  


-12'd172,  12'd9,  12'd7,  -12'd340,  12'd10,  -12'd92,  
-12'd22,  -12'd213,  -12'd355,  -12'd400,  -12'd482,  -12'd360,  
12'd122,  -12'd149,  -12'd0,  -12'd240,  12'd319,  12'd64,  
-12'd211,  -12'd81,  -12'd338,  12'd87,  12'd68,  -12'd36,  
12'd269,  12'd24,  12'd108,  12'd106,  12'd207,  12'd370,  
-12'd109,  -12'd107,  -12'd246,  -12'd186,  -12'd74,  -12'd90,  
12'd56,  12'd10,  -12'd196,  -12'd84,  -12'd59,  -12'd153,  
12'd315,  12'd388,  -12'd163,  12'd216,  -12'd257,  -12'd282,  
-12'd164,  12'd22,  -12'd325,  -12'd289,  12'd93,  -12'd652,  
-12'd271,  -12'd209,  -12'd392,  -12'd523,  -12'd215,  12'd6,  
12'd20,  12'd348,  -12'd224,  12'd246,  12'd133,  -12'd248,  
-12'd119,  -12'd415,  -12'd107,  -12'd403,  12'd112,  12'd398,  
-12'd3,  12'd52,  -12'd76,  -12'd283,  -12'd262,  -12'd10,  
-12'd103,  12'd143,  12'd430,  12'd163,  12'd59,  12'd262,  
-12'd213,  -12'd226,  -12'd164,  12'd15,  -12'd288,  -12'd45,  
-12'd60,  -12'd259,  12'd287,  12'd131,  12'd248,  12'd157,  

12'd52,  12'd57,  -12'd191,  -12'd205,  -12'd335,  -12'd421,  
-12'd81,  12'd178,  12'd152,  12'd126,  -12'd341,  -12'd144,  
-12'd241,  -12'd214,  -12'd468,  -12'd94,  12'd30,  -12'd663,  
12'd117,  12'd133,  12'd195,  12'd187,  -12'd91,  12'd104,  
12'd174,  -12'd175,  12'd369,  -12'd108,  12'd226,  12'd189,  
12'd178,  -12'd69,  12'd25,  12'd273,  -12'd370,  12'd94,  
-12'd32,  12'd92,  12'd491,  12'd79,  -12'd192,  -12'd47,  
12'd39,  -12'd265,  12'd100,  12'd187,  -12'd369,  -12'd165,  
12'd225,  12'd176,  12'd27,  -12'd257,  12'd51,  12'd176,  
-12'd123,  -12'd92,  -12'd449,  -12'd172,  -12'd250,  -12'd730,  
12'd123,  12'd11,  12'd22,  12'd113,  12'd156,  -12'd298,  
12'd68,  -12'd22,  12'd96,  -12'd10,  -12'd77,  12'd261,  
-12'd153,  12'd302,  12'd310,  12'd40,  12'd12,  12'd225,  
12'd20,  -12'd135,  12'd240,  -12'd295,  12'd69,  12'd245,  
-12'd199,  12'd58,  12'd21,  12'd36,  -12'd114,  -12'd165,  
12'd350,  12'd338,  12'd101,  12'd26,  12'd472,  -12'd322,  

12'd142,  12'd454,  -12'd163,  12'd120,  -12'd110,  -12'd531,  
12'd202,  -12'd38,  12'd56,  12'd138,  -12'd369,  -12'd60,  
-12'd321,  12'd254,  -12'd0,  12'd22,  -12'd473,  -12'd356,  
12'd345,  12'd54,  -12'd11,  12'd258,  -12'd149,  -12'd112,  
-12'd66,  12'd21,  12'd82,  -12'd417,  12'd308,  12'd347,  
12'd265,  12'd32,  12'd278,  12'd48,  12'd87,  -12'd376,  
12'd34,  12'd46,  12'd138,  -12'd24,  12'd7,  12'd231,  
12'd35,  -12'd59,  12'd401,  12'd133,  -12'd754,  12'd3,  
-12'd55,  12'd66,  12'd214,  -12'd5,  12'd386,  12'd249,  
-12'd354,  12'd71,  -12'd142,  -12'd44,  12'd426,  12'd360,  
12'd233,  12'd42,  12'd47,  12'd290,  12'd259,  -12'd248,  
12'd127,  12'd214,  -12'd344,  -12'd252,  12'd311,  12'd249,  
-12'd309,  12'd245,  -12'd31,  12'd208,  12'd157,  12'd106,  
-12'd147,  -12'd234,  -12'd324,  -12'd265,  -12'd203,  -12'd199,  
-12'd39,  12'd332,  -12'd91,  12'd250,  -12'd321,  12'd43,  
12'd364,  12'd123,  12'd259,  12'd309,  12'd681,  -12'd181,  

-12'd16,  -12'd65,  12'd386,  -12'd55,  -12'd155,  12'd200,  
12'd509,  12'd203,  12'd85,  12'd165,  -12'd253,  12'd441,  
12'd420,  12'd507,  12'd35,  12'd37,  -12'd201,  12'd488,  
12'd51,  12'd358,  12'd37,  12'd103,  -12'd202,  12'd323,  
-12'd130,  -12'd250,  12'd115,  -12'd223,  -12'd13,  12'd179,  
12'd302,  -12'd81,  -12'd250,  12'd262,  12'd31,  -12'd88,  
-12'd88,  12'd55,  12'd286,  -12'd227,  -12'd371,  12'd254,  
12'd32,  -12'd246,  12'd137,  12'd220,  -12'd410,  12'd232,  
-12'd158,  12'd325,  -12'd233,  12'd181,  12'd221,  -12'd408,  
-12'd185,  12'd305,  12'd255,  12'd26,  -12'd146,  12'd334,  
12'd392,  12'd160,  12'd181,  12'd47,  12'd607,  -12'd20,  
12'd14,  12'd109,  -12'd70,  12'd179,  -12'd90,  -12'd273,  
12'd167,  -12'd196,  12'd241,  -12'd297,  -12'd16,  -12'd102,  
12'd110,  -12'd11,  12'd72,  -12'd238,  -12'd488,  12'd10,  
-12'd15,  -12'd90,  -12'd43,  12'd16,  -12'd299,  -12'd49,  
-12'd96,  12'd162,  -12'd139,  12'd353,  12'd320,  12'd23,  

12'd122,  -12'd252,  12'd485,  12'd318,  -12'd284,  12'd407,  
12'd178,  -12'd256,  12'd58,  -12'd30,  12'd154,  12'd250,  
12'd227,  -12'd423,  12'd38,  12'd138,  -12'd368,  12'd296,  
-12'd36,  -12'd181,  12'd82,  12'd94,  -12'd83,  12'd234,  
12'd111,  -12'd213,  -12'd275,  12'd266,  -12'd723,  -12'd479,  
12'd14,  -12'd54,  12'd243,  12'd35,  -12'd154,  12'd304,  
-12'd217,  -12'd216,  -12'd244,  -12'd202,  -12'd722,  12'd76,  
12'd37,  12'd296,  12'd163,  12'd68,  -12'd38,  -12'd82,  
-12'd128,  -12'd69,  12'd176,  12'd37,  12'd319,  12'd38,  
-12'd84,  -12'd105,  12'd198,  12'd221,  12'd50,  12'd323,  
12'd114,  12'd430,  12'd448,  -12'd203,  12'd325,  12'd363,  
12'd345,  -12'd331,  12'd4,  -12'd5,  -12'd409,  -12'd57,  
-12'd131,  -12'd162,  -12'd18,  12'd201,  12'd34,  12'd195,  
12'd187,  12'd62,  12'd87,  12'd209,  -12'd653,  12'd223,  
12'd17,  12'd185,  12'd97,  12'd96,  12'd91,  12'd90,  
12'd153,  -12'd581,  -12'd91,  12'd153,  -12'd17,  -12'd328,  


-12'd86,  -12'd318,  -12'd299,  12'd146,  12'd36,  -12'd627,  
12'd135,  -12'd88,  12'd48,  12'd157,  -12'd128,  -12'd457,  
12'd43,  12'd245,  -12'd23,  12'd444,  12'd353,  -12'd489,  
-12'd108,  12'd11,  -12'd341,  12'd40,  -12'd320,  -12'd337,  
12'd133,  -12'd107,  -12'd55,  12'd339,  12'd225,  12'd414,  
12'd455,  12'd147,  -12'd225,  -12'd41,  12'd370,  -12'd163,  
-12'd295,  12'd323,  12'd211,  12'd95,  12'd37,  -12'd237,  
-12'd351,  -12'd23,  12'd187,  12'd208,  -12'd7,  12'd108,  
12'd200,  12'd492,  -12'd433,  -12'd146,  -12'd48,  -12'd40,  
-12'd167,  12'd78,  -12'd12,  -12'd297,  12'd382,  -12'd106,  
12'd152,  -12'd146,  12'd3,  12'd349,  -12'd422,  -12'd183,  
12'd264,  -12'd32,  12'd23,  12'd215,  12'd464,  12'd139,  
12'd1,  12'd418,  12'd366,  12'd268,  12'd156,  12'd132,  
12'd56,  12'd225,  12'd51,  12'd390,  -12'd47,  12'd346,  
-12'd262,  -12'd413,  12'd73,  12'd152,  -12'd706,  12'd281,  
12'd30,  -12'd13,  12'd146,  12'd173,  12'd65,  12'd302,  

-12'd31,  12'd280,  12'd74,  12'd49,  12'd256,  -12'd406,  
-12'd323,  12'd75,  12'd423,  -12'd219,  -12'd22,  12'd600,  
-12'd548,  -12'd47,  -12'd65,  -12'd210,  -12'd172,  -12'd62,  
12'd241,  12'd66,  -12'd50,  12'd555,  -12'd32,  -12'd270,  
12'd403,  12'd42,  12'd82,  -12'd217,  12'd123,  12'd176,  
-12'd449,  -12'd79,  -12'd252,  12'd355,  12'd103,  12'd175,  
12'd98,  12'd356,  12'd318,  -12'd33,  -12'd635,  12'd329,  
12'd57,  -12'd35,  -12'd384,  12'd461,  -12'd162,  -12'd203,  
-12'd253,  -12'd8,  12'd342,  -12'd415,  -12'd152,  -12'd16,  
-12'd31,  12'd193,  12'd296,  -12'd80,  12'd515,  -12'd207,  
-12'd11,  -12'd13,  -12'd162,  12'd180,  -12'd166,  -12'd12,  
12'd135,  12'd220,  -12'd243,  12'd73,  12'd310,  12'd97,  
-12'd141,  -12'd174,  12'd206,  12'd429,  12'd71,  12'd192,  
12'd103,  12'd131,  12'd143,  -12'd325,  12'd260,  12'd220,  
-12'd259,  12'd168,  -12'd338,  12'd111,  -12'd348,  -12'd211,  
12'd217,  -12'd127,  12'd91,  -12'd267,  12'd86,  12'd303,  

-12'd162,  12'd161,  12'd89,  12'd56,  12'd214,  -12'd33,  
-12'd312,  -12'd169,  -12'd5,  -12'd178,  -12'd13,  12'd557,  
-12'd252,  12'd113,  -12'd138,  12'd109,  -12'd276,  -12'd197,  
12'd298,  12'd17,  12'd208,  12'd241,  12'd129,  -12'd588,  
12'd310,  -12'd289,  -12'd152,  12'd125,  12'd67,  12'd100,  
-12'd392,  12'd62,  12'd135,  12'd276,  -12'd199,  -12'd343,  
12'd230,  -12'd221,  12'd541,  12'd64,  -12'd370,  12'd233,  
12'd213,  12'd6,  -12'd266,  12'd316,  -12'd346,  -12'd140,  
-12'd65,  -12'd319,  -12'd200,  -12'd173,  -12'd316,  12'd137,  
12'd7,  -12'd5,  12'd129,  -12'd7,  12'd268,  -12'd58,  
12'd156,  12'd215,  -12'd241,  12'd261,  12'd198,  12'd173,  
12'd219,  12'd118,  -12'd133,  -12'd9,  -12'd248,  12'd195,  
12'd316,  12'd207,  -12'd120,  12'd343,  12'd58,  12'd33,  
-12'd340,  12'd48,  -12'd283,  -12'd53,  -12'd499,  -12'd326,  
12'd263,  12'd592,  12'd87,  12'd149,  -12'd621,  12'd149,  
12'd157,  -12'd405,  12'd140,  12'd47,  12'd8,  12'd290,  

-12'd574,  12'd530,  12'd516,  12'd248,  -12'd333,  12'd556,  
12'd52,  -12'd225,  -12'd228,  -12'd66,  -12'd520,  12'd148,  
12'd34,  12'd282,  12'd261,  12'd554,  -12'd658,  12'd145,  
12'd301,  12'd208,  12'd69,  12'd404,  12'd473,  -12'd307,  
-12'd263,  12'd46,  -12'd238,  -12'd395,  12'd354,  12'd406,  
12'd379,  12'd379,  12'd153,  12'd224,  -12'd194,  -12'd514,  
12'd69,  -12'd553,  -12'd92,  -12'd60,  -12'd244,  12'd186,  
12'd77,  12'd203,  12'd149,  12'd377,  12'd363,  12'd65,  
12'd226,  -12'd64,  -12'd231,  -12'd33,  12'd402,  12'd27,  
12'd343,  -12'd236,  -12'd315,  12'd349,  12'd30,  -12'd637,  
12'd246,  -12'd358,  12'd207,  12'd97,  12'd216,  12'd398,  
12'd129,  12'd41,  12'd285,  -12'd163,  -12'd245,  12'd205,  
12'd442,  12'd92,  12'd130,  12'd409,  12'd57,  -12'd176,  
-12'd450,  12'd80,  -12'd111,  12'd274,  -12'd596,  12'd472,  
12'd436,  12'd20,  12'd378,  -12'd49,  -12'd7,  -12'd421,  
12'd284,  -12'd167,  12'd150,  -12'd188,  -12'd283,  -12'd528,  

12'd383,  -12'd133,  12'd196,  12'd72,  -12'd793,  12'd650,  
12'd1,  -12'd32,  -12'd264,  12'd103,  -12'd199,  12'd225,  
12'd220,  12'd36,  -12'd220,  -12'd35,  -12'd530,  12'd15,  
12'd312,  12'd433,  12'd271,  12'd69,  12'd398,  12'd95,  
-12'd132,  -12'd97,  -12'd24,  -12'd269,  12'd135,  12'd311,  
12'd217,  12'd192,  -12'd107,  12'd447,  -12'd299,  12'd30,  
12'd120,  12'd152,  -12'd592,  -12'd353,  -12'd564,  -12'd472,  
12'd105,  12'd329,  -12'd265,  12'd450,  12'd185,  12'd86,  
12'd294,  12'd290,  -12'd249,  12'd188,  12'd285,  12'd96,  
12'd513,  -12'd159,  -12'd21,  12'd130,  12'd271,  -12'd280,  
12'd21,  -12'd281,  12'd136,  -12'd264,  -12'd734,  12'd304,  
-12'd242,  12'd237,  12'd685,  -12'd384,  -12'd200,  12'd878,  
12'd51,  12'd181,  12'd292,  12'd75,  12'd207,  12'd135,  
-12'd47,  12'd277,  12'd146,  12'd426,  -12'd585,  12'd233,  
-12'd26,  12'd86,  12'd7,  12'd5,  12'd45,  -12'd329,  
12'd436,  -12'd53,  12'd85,  -12'd159,  -12'd334,  12'd174,  


12'd250,  12'd235,  12'd33,  -12'd72,  12'd432,  -12'd232,  
-12'd47,  12'd177,  12'd238,  -12'd192,  -12'd22,  12'd295,  
12'd305,  12'd367,  12'd211,  12'd177,  12'd311,  -12'd419,  
12'd53,  12'd142,  12'd243,  12'd397,  12'd171,  -12'd255,  
-12'd400,  -12'd315,  12'd88,  -12'd100,  -12'd482,  12'd46,  
12'd157,  12'd254,  -12'd171,  12'd359,  -12'd15,  12'd62,  
-12'd577,  12'd292,  12'd494,  12'd319,  -12'd372,  12'd79,  
-12'd57,  -12'd301,  12'd199,  12'd159,  -12'd341,  12'd144,  
12'd108,  12'd403,  12'd413,  12'd42,  -12'd230,  12'd654,  
12'd332,  12'd281,  -12'd340,  -12'd44,  12'd258,  12'd124,  
-12'd493,  -12'd14,  -12'd333,  12'd346,  -12'd355,  12'd217,  
-12'd36,  -12'd210,  -12'd257,  12'd6,  12'd201,  12'd172,  
-12'd92,  -12'd187,  12'd23,  12'd331,  12'd131,  12'd239,  
-12'd60,  12'd33,  -12'd134,  -12'd83,  -12'd56,  12'd49,  
12'd214,  -12'd321,  12'd99,  -12'd211,  -12'd448,  -12'd29,  
12'd37,  -12'd208,  -12'd265,  -12'd166,  -12'd178,  -12'd15,  

-12'd398,  12'd406,  12'd393,  12'd54,  12'd203,  12'd418,  
-12'd290,  12'd267,  12'd666,  -12'd113,  -12'd252,  12'd335,  
12'd104,  -12'd46,  -12'd101,  -12'd27,  12'd149,  -12'd486,  
12'd100,  -12'd28,  -12'd208,  12'd133,  12'd108,  -12'd231,  
-12'd122,  -12'd40,  12'd26,  12'd12,  12'd20,  12'd29,  
-12'd483,  12'd126,  12'd163,  12'd103,  -12'd169,  12'd15,  
-12'd17,  -12'd108,  12'd196,  12'd182,  -12'd501,  -12'd36,  
-12'd405,  -12'd261,  -12'd69,  -12'd15,  -12'd888,  12'd22,  
-12'd307,  12'd241,  12'd271,  -12'd230,  -12'd134,  12'd308,  
12'd9,  12'd219,  12'd179,  12'd277,  12'd315,  12'd159,  
-12'd282,  12'd60,  -12'd63,  -12'd158,  12'd69,  12'd74,  
-12'd74,  12'd131,  12'd59,  -12'd15,  12'd173,  12'd3,  
12'd484,  -12'd339,  -12'd140,  -12'd140,  -12'd81,  12'd35,  
12'd109,  12'd143,  12'd191,  -12'd208,  12'd112,  12'd384,  
12'd362,  12'd274,  -12'd298,  -12'd18,  -12'd325,  -12'd38,  
12'd98,  -12'd69,  12'd112,  -12'd192,  12'd100,  -12'd152,  

-12'd431,  -12'd19,  -12'd79,  12'd234,  -12'd312,  12'd219,  
12'd135,  -12'd261,  12'd170,  -12'd431,  -12'd704,  12'd232,  
-12'd363,  12'd124,  -12'd158,  12'd61,  -12'd325,  -12'd261,  
12'd254,  12'd117,  -12'd59,  12'd163,  -12'd84,  -12'd329,  
12'd282,  12'd76,  12'd390,  -12'd0,  12'd11,  -12'd25,  
-12'd457,  -12'd111,  -12'd206,  -12'd424,  -12'd181,  12'd433,  
12'd449,  -12'd209,  -12'd83,  12'd76,  -12'd585,  12'd48,  
-12'd215,  -12'd364,  -12'd180,  12'd243,  -12'd259,  -12'd373,  
12'd61,  -12'd609,  -12'd230,  -12'd261,  -12'd413,  12'd252,  
12'd242,  -12'd213,  -12'd100,  -12'd162,  -12'd66,  -12'd329,  
-12'd249,  -12'd99,  -12'd24,  12'd275,  12'd253,  -12'd383,  
12'd97,  12'd147,  12'd244,  -12'd264,  12'd206,  12'd134,  
12'd216,  -12'd34,  -12'd481,  12'd360,  12'd21,  -12'd106,  
-12'd145,  -12'd234,  -12'd110,  -12'd341,  -12'd127,  -12'd88,  
12'd69,  12'd325,  12'd3,  12'd574,  -12'd295,  -12'd244,  
-12'd123,  12'd10,  -12'd278,  -12'd378,  12'd181,  -12'd455,  

12'd30,  -12'd108,  -12'd344,  12'd56,  -12'd1088,  -12'd259,  
-12'd171,  -12'd181,  -12'd382,  -12'd85,  -12'd772,  -12'd173,  
-12'd267,  12'd2,  12'd202,  12'd205,  -12'd828,  12'd268,  
-12'd35,  -12'd186,  -12'd267,  12'd358,  12'd294,  -12'd136,  
12'd179,  12'd372,  -12'd122,  12'd35,  12'd429,  -12'd494,  
12'd231,  -12'd282,  -12'd189,  12'd183,  -12'd660,  -12'd160,  
12'd68,  -12'd213,  -12'd538,  -12'd373,  -12'd171,  -12'd445,  
12'd385,  -12'd61,  -12'd262,  12'd78,  -12'd153,  -12'd603,  
12'd564,  12'd310,  -12'd231,  -12'd285,  -12'd101,  -12'd250,  
-12'd37,  12'd51,  -12'd90,  -12'd38,  12'd121,  -12'd489,  
-12'd187,  -12'd656,  -12'd465,  -12'd239,  -12'd24,  -12'd226,  
-12'd261,  -12'd98,  12'd229,  12'd320,  -12'd213,  12'd257,  
-12'd110,  -12'd219,  -12'd238,  12'd436,  12'd244,  -12'd558,  
-12'd244,  12'd20,  12'd95,  12'd16,  -12'd569,  12'd321,  
12'd216,  12'd112,  -12'd115,  12'd371,  12'd162,  -12'd94,  
-12'd330,  12'd113,  -12'd37,  -12'd89,  -12'd159,  12'd101,  

-12'd90,  12'd45,  -12'd57,  12'd139,  -12'd369,  12'd128,  
12'd129,  12'd371,  12'd94,  12'd39,  -12'd375,  12'd488,  
12'd265,  -12'd48,  12'd129,  12'd124,  -12'd228,  -12'd300,  
12'd545,  12'd125,  12'd24,  12'd99,  12'd256,  -12'd130,  
12'd135,  12'd80,  12'd72,  -12'd63,  12'd119,  -12'd141,  
12'd298,  -12'd25,  12'd120,  12'd498,  -12'd30,  -12'd486,  
-12'd22,  12'd271,  -12'd124,  -12'd339,  -12'd43,  -12'd24,  
12'd385,  12'd98,  -12'd73,  12'd255,  12'd385,  -12'd536,  
12'd621,  -12'd201,  -12'd466,  -12'd77,  12'd553,  -12'd16,  
12'd84,  -12'd13,  -12'd275,  12'd163,  -12'd395,  -12'd364,  
-12'd279,  -12'd229,  -12'd650,  -12'd550,  12'd127,  -12'd311,  
-12'd304,  12'd34,  -12'd41,  12'd143,  -12'd832,  12'd628,  
12'd56,  -12'd47,  -12'd32,  -12'd250,  12'd333,  -12'd168,  
12'd329,  -12'd156,  12'd384,  12'd326,  -12'd467,  12'd69,  
12'd374,  12'd17,  12'd38,  12'd342,  -12'd16,  -12'd30,  
12'd6,  -12'd177,  12'd93,  12'd180,  -12'd359,  12'd454,  


-12'd125,  12'd12,  -12'd167,  -12'd475,  12'd278,  12'd473,  
-12'd456,  12'd180,  -12'd52,  -12'd44,  -12'd136,  -12'd32,  
12'd538,  -12'd178,  -12'd189,  12'd101,  -12'd66,  -12'd152,  
-12'd355,  -12'd317,  12'd104,  -12'd39,  -12'd188,  -12'd138,  
12'd168,  12'd141,  -12'd105,  -12'd360,  12'd40,  -12'd161,  
-12'd374,  12'd390,  12'd220,  -12'd86,  -12'd277,  12'd230,  
-12'd57,  12'd338,  12'd552,  12'd81,  -12'd304,  12'd17,  
-12'd235,  -12'd387,  12'd227,  12'd67,  12'd220,  -12'd493,  
-12'd353,  12'd664,  12'd757,  12'd428,  -12'd769,  12'd447,  
12'd385,  -12'd227,  12'd139,  12'd101,  -12'd152,  12'd24,  
-12'd290,  12'd193,  12'd82,  -12'd65,  -12'd156,  12'd283,  
-12'd330,  12'd143,  -12'd359,  -12'd77,  -12'd341,  12'd106,  
12'd113,  -12'd251,  -12'd550,  -12'd412,  12'd176,  -12'd139,  
-12'd68,  12'd319,  12'd286,  12'd132,  -12'd292,  -12'd36,  
-12'd61,  -12'd114,  -12'd170,  -12'd55,  -12'd410,  -12'd76,  
12'd78,  -12'd124,  -12'd325,  -12'd306,  12'd352,  -12'd5,  

-12'd280,  12'd98,  12'd282,  -12'd125,  -12'd416,  12'd169,  
-12'd353,  12'd252,  12'd193,  -12'd87,  -12'd717,  12'd392,  
12'd109,  12'd179,  12'd202,  -12'd28,  12'd92,  -12'd405,  
-12'd157,  -12'd534,  -12'd115,  12'd89,  -12'd492,  12'd242,  
-12'd77,  -12'd59,  -12'd32,  -12'd265,  12'd12,  12'd476,  
-12'd87,  12'd57,  12'd17,  -12'd64,  -12'd166,  12'd271,  
12'd279,  12'd159,  -12'd23,  12'd91,  -12'd577,  12'd409,  
-12'd482,  -12'd73,  -12'd407,  -12'd211,  -12'd227,  -12'd8,  
12'd300,  12'd312,  12'd462,  12'd288,  -12'd732,  12'd543,  
12'd429,  12'd59,  -12'd271,  12'd266,  12'd243,  -12'd583,  
12'd96,  -12'd500,  -12'd392,  -12'd271,  12'd509,  -12'd43,  
-12'd17,  12'd202,  12'd43,  -12'd121,  -12'd143,  -12'd13,  
-12'd13,  -12'd382,  -12'd193,  -12'd154,  12'd556,  -12'd173,  
-12'd175,  -12'd69,  12'd429,  12'd49,  -12'd157,  -12'd29,  
-12'd315,  12'd67,  -12'd115,  -12'd518,  -12'd231,  -12'd201,  
12'd242,  12'd84,  -12'd109,  -12'd35,  12'd390,  -12'd207,  

-12'd273,  12'd236,  -12'd123,  12'd263,  -12'd789,  12'd46,  
12'd432,  -12'd419,  -12'd196,  12'd76,  -12'd199,  12'd76,  
-12'd125,  12'd330,  -12'd233,  12'd22,  -12'd244,  12'd123,  
-12'd231,  -12'd478,  -12'd266,  12'd192,  -12'd202,  -12'd247,  
-12'd311,  12'd193,  12'd156,  -12'd21,  -12'd106,  12'd67,  
-12'd210,  -12'd606,  12'd83,  -12'd117,  -12'd295,  12'd75,  
12'd157,  -12'd372,  -12'd143,  -12'd30,  -12'd280,  -12'd267,  
-12'd219,  -12'd229,  12'd175,  -12'd118,  -12'd7,  -12'd113,  
12'd341,  12'd174,  -12'd190,  12'd110,  -12'd80,  -12'd134,  
12'd224,  12'd339,  -12'd303,  -12'd137,  12'd100,  -12'd540,  
-12'd355,  12'd72,  -12'd565,  -12'd298,  12'd110,  -12'd794,  
-12'd392,  12'd7,  12'd153,  12'd254,  -12'd236,  12'd485,  
-12'd195,  12'd44,  -12'd243,  -12'd175,  12'd300,  -12'd33,  
-12'd122,  12'd62,  12'd200,  -12'd171,  12'd304,  -12'd187,  
-12'd106,  -12'd283,  -12'd140,  12'd33,  -12'd387,  -12'd434,  
-12'd65,  12'd135,  -12'd115,  -12'd324,  12'd250,  12'd488,  

12'd359,  -12'd240,  -12'd304,  12'd165,  -12'd437,  -12'd213,  
-12'd44,  12'd22,  12'd208,  -12'd157,  -12'd155,  12'd185,  
12'd77,  12'd98,  12'd145,  12'd100,  -12'd462,  12'd497,  
-12'd391,  -12'd499,  -12'd436,  -12'd101,  -12'd442,  -12'd423,  
12'd131,  12'd7,  12'd297,  -12'd59,  -12'd77,  -12'd114,  
12'd47,  -12'd33,  -12'd177,  -12'd43,  -12'd65,  -12'd421,  
12'd11,  12'd150,  -12'd246,  12'd92,  12'd389,  -12'd376,  
-12'd317,  -12'd291,  12'd47,  -12'd255,  -12'd114,  12'd86,  
-12'd372,  -12'd42,  -12'd304,  -12'd482,  12'd43,  12'd117,  
12'd183,  12'd293,  -12'd155,  12'd30,  12'd637,  12'd101,  
-12'd262,  -12'd313,  -12'd403,  -12'd617,  12'd183,  -12'd441,  
12'd86,  -12'd501,  -12'd125,  12'd105,  12'd34,  12'd116,  
-12'd612,  -12'd180,  -12'd8,  -12'd464,  -12'd47,  -12'd204,  
12'd119,  12'd309,  12'd368,  -12'd6,  -12'd309,  12'd40,  
12'd272,  12'd19,  -12'd240,  12'd119,  -12'd206,  -12'd53,  
-12'd433,  12'd91,  12'd251,  -12'd96,  -12'd154,  12'd4,  

-12'd72,  -12'd244,  -12'd489,  12'd231,  -12'd223,  -12'd360,  
-12'd205,  -12'd14,  12'd455,  12'd206,  -12'd290,  12'd473,  
12'd346,  -12'd362,  -12'd266,  12'd372,  -12'd136,  12'd31,  
-12'd100,  -12'd232,  -12'd98,  -12'd206,  -12'd232,  -12'd439,  
12'd112,  -12'd63,  -12'd88,  12'd38,  -12'd41,  -12'd29,  
-12'd41,  -12'd406,  -12'd243,  -12'd141,  -12'd456,  -12'd94,  
12'd187,  12'd494,  -12'd75,  -12'd50,  12'd158,  12'd143,  
-12'd351,  -12'd216,  -12'd253,  -12'd138,  -12'd31,  12'd173,  
12'd244,  -12'd477,  -12'd147,  -12'd132,  12'd9,  -12'd49,  
-12'd2,  -12'd248,  12'd150,  -12'd249,  12'd101,  -12'd402,  
-12'd403,  12'd428,  -12'd108,  -12'd336,  12'd137,  -12'd277,  
-12'd47,  -12'd23,  -12'd40,  12'd68,  12'd105,  -12'd698,  
-12'd661,  -12'd300,  12'd65,  -12'd468,  -12'd494,  12'd271,  
12'd435,  12'd322,  -12'd85,  12'd52,  -12'd349,  -12'd79,  
12'd218,  -12'd501,  12'd108,  -12'd16,  -12'd169,  -12'd144,  
-12'd91,  -12'd109,  -12'd21,  12'd213,  -12'd318,  12'd49
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
	


endmodule


module bias_fc1_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC1-1][0:`OUTPUT_NUM_FC1-1][`WD_BIAS:0] weight	 = {
-24'd219560,  -24'd253697,  -24'd55433,  -24'd97677,  24'd293697,  -24'd243881,  24'd320084,  24'd224550,  24'd239030,  24'd511222,  24'd91710,  24'd236129,  24'd189478,  24'd189715,  24'd237750,  24'd85050,  
24'd84279,  -24'd41102,  24'd389770,  24'd141391,  -24'd114359,  24'd179309,  24'd335280,  24'd91496,  -24'd304524,  24'd51767,  24'd50531,  24'd398249,  24'd125193,  24'd59246,  24'd302096,  -24'd391546,  
-24'd8719,  -24'd143200,  24'd86710,  -24'd121286,  -24'd17574,  24'd193986,  24'd334251,  24'd418338,  -24'd29725,  -24'd164781,  24'd19566,  24'd369659,  24'd369117,  24'd485986,  24'd255667,  24'd184972,  
-24'd350874,  24'd83616,  -24'd113753,  24'd50318,  -24'd218172,  24'd245365,  -24'd212866,  -24'd167942,  24'd24266,  -24'd290894,  -24'd45370,  24'd333035,  24'd76391,  24'd331919,  24'd249570,  24'd116175,  
24'd314113,  24'd322302,  -24'd387295,  -24'd139803,  24'd555959,  24'd41557,  -24'd71756,  24'd250106,  24'd125286,  24'd209370,  -24'd167080,  24'd330490,  24'd186924,  24'd87729,  -24'd220844,  24'd340936,  
-24'd135930,  24'd117423,  24'd224274,  -24'd3834,  -24'd49645,  -24'd105418,  24'd52762,  24'd96732,  -24'd152523,  24'd141711,  24'd257837,  -24'd91013,  24'd178395,  24'd55568,  -24'd93767,  -24'd131308,  
24'd155983,  -24'd449369,  24'd184192,  -24'd39257,  -24'd140313,  24'd360847,  24'd255272,  24'd73788,  -24'd213748,  24'd163158,  24'd149546,  24'd206663,  -24'd58642,  -24'd77157,  -24'd41775,  24'd140758,  
24'd396969,  24'd190957,  24'd87027,  -24'd48891,  24'd157309,  -24'd282668,  -24'd283377,  -24'd195665
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule

module wieght_fc1_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1*`OUTPUT_BATCH_FC1)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_CONV2*`OUTPUT_NUM_FC1 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC1*`KERNEL_SIZE_FC1*`KERNEL_SIZE_FC1-1][0:`OUTPUT_NUM_FC1-1][0:`OUTPUT_NUM_CONV2-1][`WD:0] weight	 = {
-12'd88,  12'd49,  -12'd52,  12'd500,  -12'd4,  12'd0,  12'd120,  -12'd438,  12'd224,  12'd139,  -12'd70,  -12'd133,  12'd205,  -12'd230,  -12'd178,  -12'd48,  
12'd439,  12'd46,  12'd240,  12'd211,  -12'd217,  12'd165,  -12'd288,  12'd245,  12'd42,  -12'd29,  12'd4,  12'd65,  12'd252,  -12'd140,  -12'd13,  12'd76,  
12'd161,  -12'd278,  12'd85,  -12'd252,  -12'd338,  -12'd155,  12'd42,  -12'd287,  12'd121,  -12'd235,  12'd429,  12'd256,  12'd315,  -12'd146,  -12'd220,  12'd495,  
12'd120,  12'd53,  12'd183,  12'd0,  -12'd200,  12'd334,  12'd429,  12'd143,  12'd321,  -12'd8,  12'd285,  12'd3,  12'd175,  12'd352,  -12'd111,  -12'd43,  
12'd458,  12'd409,  -12'd328,  12'd160,  12'd469,  12'd336,  12'd324,  12'd289,  12'd195,  -12'd130,  12'd46,  12'd329,  12'd457,  12'd175,  -12'd508,  12'd132,  
12'd257,  12'd170,  -12'd254,  12'd186,  12'd211,  -12'd85,  12'd193,  -12'd403,  -12'd139,  -12'd200,  12'd526,  -12'd116,  -12'd34,  -12'd229,  12'd382,  -12'd13,  
12'd40,  12'd133,  -12'd148,  -12'd168,  -12'd36,  12'd196,  12'd97,  -12'd14,  12'd146,  12'd91,  12'd432,  12'd121,  -12'd288,  -12'd151,  -12'd475,  -12'd355,  
12'd83,  -12'd266,  -12'd140,  -12'd223,  -12'd25,  12'd106,  12'd51,  -12'd248,  12'd68,  12'd349,  -12'd50,  12'd119,  12'd417,  -12'd48,  -12'd184,  12'd149,  
12'd281,  -12'd335,  -12'd240,  -12'd333,  -12'd21,  12'd63,  -12'd157,  -12'd308,  -12'd287,  -12'd441,  -12'd188,  -12'd170,  12'd265,  12'd358,  12'd148,  12'd111,  
-12'd89,  -12'd36,  -12'd752,  -12'd148,  -12'd208,  -12'd111,  -12'd23,  -12'd50,  -12'd267,  -12'd301,  12'd174,  -12'd213,  -12'd182,  -12'd186,  12'd186,  -12'd322,  
-12'd92,  12'd35,  12'd411,  -12'd440,  -12'd111,  -12'd253,  -12'd49,  -12'd239,  -12'd121,  -12'd260,  -12'd307,  12'd138,  12'd161,  -12'd56,  -12'd13,  -12'd40,  
-12'd25,  12'd337,  12'd221,  -12'd353,  -12'd283,  12'd6,  12'd217,  -12'd96,  12'd147,  12'd126,  -12'd328,  -12'd62,  -12'd304,  12'd360,  -12'd261,  -12'd109,  
-12'd2,  -12'd164,  -12'd224,  -12'd304,  -12'd205,  -12'd267,  -12'd285,  -12'd358,  -12'd303,  -12'd175,  -12'd475,  -12'd205,  12'd88,  12'd382,  -12'd171,  -12'd133,  
12'd4,  -12'd163,  12'd307,  12'd196,  -12'd3,  -12'd658,  -12'd115,  -12'd114,  12'd19,  12'd230,  -12'd370,  -12'd234,  12'd18,  12'd236,  -12'd271,  -12'd6,  
-12'd543,  -12'd343,  12'd140,  12'd175,  -12'd60,  -12'd467,  12'd38,  -12'd380,  -12'd3,  12'd395,  -12'd28,  12'd201,  -12'd254,  -12'd112,  -12'd5,  -12'd499,  
-12'd125,  -12'd166,  12'd67,  12'd336,  12'd238,  -12'd34,  -12'd577,  -12'd74,  12'd168,  -12'd7,  -12'd320,  -12'd314,  12'd102,  -12'd15,  12'd452,  -12'd61,  
-12'd216,  -12'd366,  -12'd72,  12'd601,  12'd197,  -12'd51,  -12'd162,  12'd186,  -12'd193,  -12'd14,  12'd416,  -12'd276,  -12'd39,  -12'd117,  -12'd66,  -12'd345,  
12'd18,  -12'd52,  12'd111,  12'd46,  -12'd93,  -12'd400,  -12'd682,  12'd38,  -12'd605,  12'd342,  -12'd55,  -12'd197,  12'd196,  12'd2,  -12'd85,  12'd340,  
-12'd61,  -12'd243,  12'd116,  12'd183,  -12'd354,  12'd38,  12'd49,  -12'd15,  -12'd168,  -12'd334,  -12'd311,  12'd343,  12'd328,  -12'd5,  12'd67,  12'd225,  
-12'd170,  -12'd235,  -12'd188,  -12'd141,  -12'd96,  -12'd56,  12'd291,  12'd76,  12'd278,  -12'd242,  12'd35,  12'd405,  -12'd80,  -12'd74,  -12'd8,  -12'd137,  
-12'd261,  12'd367,  -12'd276,  -12'd206,  12'd54,  12'd144,  -12'd267,  12'd181,  12'd689,  12'd93,  12'd544,  -12'd399,  -12'd12,  -12'd333,  12'd33,  -12'd7,  
-12'd210,  12'd77,  -12'd518,  -12'd192,  -12'd148,  -12'd208,  -12'd581,  -12'd333,  12'd313,  -12'd371,  12'd196,  12'd22,  -12'd56,  -12'd578,  12'd26,  12'd290,  
12'd34,  -12'd50,  -12'd366,  12'd45,  -12'd580,  -12'd278,  -12'd436,  12'd175,  -12'd169,  -12'd120,  12'd215,  -12'd61,  -12'd117,  12'd400,  12'd76,  -12'd30,  
-12'd218,  12'd35,  12'd491,  -12'd325,  -12'd368,  -12'd8,  12'd372,  -12'd220,  12'd9,  -12'd90,  -12'd190,  12'd84,  12'd80,  12'd586,  12'd411,  12'd205,  
12'd332,  12'd114,  12'd328,  12'd238,  -12'd2,  12'd163,  12'd336,  12'd65,  12'd60,  -12'd561,  -12'd174,  12'd210,  -12'd124,  -12'd118,  12'd230,  12'd246,  

-12'd106,  -12'd1,  -12'd66,  12'd120,  -12'd138,  12'd201,  -12'd277,  -12'd51,  -12'd381,  -12'd87,  12'd25,  12'd144,  -12'd43,  -12'd103,  12'd103,  12'd187,  
-12'd312,  -12'd341,  -12'd188,  -12'd206,  -12'd306,  -12'd232,  -12'd27,  -12'd54,  12'd28,  -12'd252,  12'd82,  12'd266,  12'd277,  12'd101,  -12'd436,  -12'd211,  
-12'd114,  -12'd209,  -12'd123,  -12'd173,  -12'd56,  12'd270,  -12'd118,  12'd171,  12'd108,  -12'd318,  -12'd105,  -12'd192,  -12'd55,  12'd91,  12'd122,  -12'd230,  
12'd137,  12'd187,  -12'd36,  12'd97,  -12'd128,  -12'd29,  -12'd425,  -12'd158,  -12'd231,  -12'd78,  -12'd445,  -12'd56,  -12'd164,  -12'd127,  12'd5,  12'd7,  
12'd351,  -12'd138,  -12'd85,  -12'd227,  12'd132,  -12'd426,  -12'd152,  -12'd86,  -12'd178,  12'd111,  -12'd414,  -12'd19,  12'd84,  12'd69,  -12'd33,  -12'd389,  
12'd63,  12'd11,  12'd274,  -12'd205,  12'd88,  12'd186,  -12'd157,  -12'd239,  -12'd113,  12'd239,  -12'd274,  12'd101,  12'd353,  12'd34,  -12'd132,  -12'd387,  
-12'd55,  -12'd100,  -12'd250,  -12'd78,  -12'd63,  -12'd89,  12'd118,  -12'd176,  -12'd263,  12'd267,  12'd160,  -12'd328,  -12'd10,  12'd122,  -12'd67,  -12'd268,  
12'd236,  -12'd212,  12'd84,  12'd187,  12'd205,  12'd190,  -12'd272,  12'd79,  12'd107,  12'd72,  -12'd70,  12'd155,  -12'd94,  -12'd71,  12'd186,  12'd170,  
-12'd10,  -12'd302,  12'd9,  -12'd234,  -12'd88,  12'd80,  12'd191,  -12'd230,  12'd49,  -12'd40,  -12'd35,  -12'd266,  -12'd496,  -12'd195,  12'd11,  -12'd459,  
12'd52,  -12'd67,  -12'd72,  -12'd198,  12'd92,  12'd31,  -12'd225,  -12'd69,  12'd78,  12'd60,  -12'd9,  -12'd49,  12'd23,  -12'd85,  -12'd389,  -12'd295,  
-12'd129,  -12'd127,  -12'd16,  -12'd394,  -12'd364,  -12'd91,  -12'd266,  -12'd4,  -12'd401,  12'd64,  12'd71,  -12'd151,  -12'd209,  12'd9,  -12'd78,  -12'd18,  
-12'd407,  -12'd379,  -12'd18,  -12'd140,  12'd156,  -12'd275,  12'd35,  -12'd62,  12'd107,  12'd288,  12'd51,  -12'd199,  12'd108,  -12'd73,  -12'd17,  12'd38,  
12'd52,  12'd22,  -12'd362,  12'd187,  12'd170,  -12'd272,  12'd31,  -12'd199,  12'd142,  -12'd169,  12'd128,  12'd275,  12'd114,  -12'd221,  12'd126,  -12'd233,  
-12'd43,  -12'd72,  -12'd186,  12'd274,  -12'd319,  12'd229,  12'd99,  -12'd114,  -12'd127,  -12'd409,  -12'd235,  -12'd206,  12'd84,  12'd129,  -12'd193,  12'd68,  
-12'd98,  -12'd67,  12'd46,  -12'd204,  12'd190,  -12'd74,  -12'd340,  12'd149,  -12'd94,  -12'd58,  -12'd139,  -12'd146,  -12'd124,  -12'd159,  -12'd235,  -12'd129,  
12'd295,  12'd94,  -12'd211,  -12'd210,  -12'd196,  -12'd120,  -12'd378,  -12'd235,  12'd201,  -12'd213,  -12'd335,  12'd22,  -12'd25,  -12'd152,  -12'd171,  -12'd191,  
-12'd404,  12'd134,  -12'd29,  12'd130,  -12'd188,  12'd95,  12'd87,  -12'd56,  -12'd369,  12'd86,  -12'd147,  -12'd300,  -12'd394,  -12'd162,  -12'd266,  12'd261,  
12'd67,  12'd241,  12'd10,  12'd188,  12'd257,  -12'd150,  12'd161,  -12'd155,  -12'd259,  12'd20,  -12'd188,  12'd247,  -12'd5,  -12'd120,  12'd113,  -12'd269,  
-12'd39,  -12'd112,  -12'd63,  -12'd160,  -12'd192,  12'd44,  -12'd254,  -12'd101,  12'd34,  12'd113,  -12'd185,  -12'd267,  -12'd350,  -12'd94,  -12'd137,  -12'd181,  
12'd55,  -12'd229,  -12'd14,  -12'd134,  -12'd247,  -12'd217,  -12'd1,  -12'd383,  -12'd25,  -12'd113,  -12'd281,  12'd181,  12'd71,  -12'd293,  12'd98,  12'd10,  
-12'd209,  12'd73,  12'd144,  -12'd245,  -12'd348,  -12'd46,  -12'd319,  12'd46,  -12'd15,  -12'd418,  12'd63,  -12'd92,  -12'd132,  -12'd424,  12'd117,  12'd24,  
12'd187,  -12'd354,  -12'd101,  -12'd77,  -12'd163,  -12'd192,  -12'd79,  12'd21,  12'd298,  -12'd79,  -12'd397,  12'd3,  12'd195,  -12'd290,  -12'd16,  -12'd238,  
12'd45,  -12'd34,  12'd331,  12'd48,  -12'd221,  -12'd97,  12'd228,  12'd62,  12'd69,  12'd241,  12'd46,  -12'd334,  -12'd157,  -12'd26,  -12'd150,  12'd198,  
-12'd179,  -12'd323,  12'd48,  -12'd294,  -12'd51,  12'd229,  -12'd83,  -12'd44,  -12'd124,  -12'd137,  -12'd39,  -12'd41,  -12'd170,  -12'd260,  12'd115,  -12'd42,  
-12'd79,  -12'd246,  12'd46,  12'd321,  -12'd132,  -12'd258,  -12'd347,  -12'd207,  12'd152,  12'd18,  12'd64,  -12'd63,  -12'd21,  -12'd231,  12'd178,  12'd131,  

-12'd217,  -12'd234,  12'd390,  -12'd216,  -12'd250,  12'd130,  -12'd618,  12'd99,  12'd310,  -12'd274,  -12'd468,  12'd60,  -12'd61,  12'd98,  12'd304,  12'd51,  
12'd62,  -12'd100,  12'd766,  -12'd93,  -12'd33,  12'd163,  12'd51,  -12'd359,  12'd66,  12'd313,  -12'd602,  12'd162,  12'd126,  -12'd104,  12'd119,  -12'd182,  
-12'd263,  12'd32,  12'd71,  -12'd300,  12'd266,  12'd85,  12'd355,  -12'd112,  -12'd129,  12'd15,  -12'd15,  12'd253,  -12'd203,  12'd965,  -12'd69,  -12'd202,  
-12'd236,  12'd241,  12'd236,  12'd222,  -12'd44,  12'd30,  12'd239,  -12'd137,  12'd332,  -12'd11,  -12'd48,  -12'd290,  -12'd313,  12'd476,  12'd133,  -12'd4,  
12'd503,  12'd619,  -12'd128,  -12'd112,  -12'd65,  -12'd66,  12'd415,  12'd163,  12'd175,  12'd47,  -12'd174,  12'd54,  -12'd180,  -12'd185,  12'd92,  12'd206,  
12'd1,  12'd48,  12'd418,  12'd325,  12'd259,  12'd106,  -12'd579,  12'd159,  -12'd336,  12'd232,  -12'd320,  -12'd49,  -12'd116,  12'd263,  -12'd4,  12'd121,  
-12'd92,  12'd247,  12'd14,  -12'd191,  -12'd50,  -12'd49,  12'd166,  12'd175,  12'd13,  12'd106,  12'd41,  -12'd17,  -12'd16,  -12'd204,  12'd134,  -12'd189,  
-12'd219,  -12'd474,  12'd237,  -12'd317,  -12'd402,  -12'd299,  12'd164,  12'd79,  12'd6,  -12'd78,  -12'd406,  -12'd230,  -12'd129,  12'd44,  12'd358,  -12'd34,  
12'd215,  12'd7,  -12'd49,  -12'd92,  -12'd300,  12'd1,  12'd17,  -12'd173,  12'd140,  -12'd271,  -12'd4,  -12'd153,  -12'd26,  12'd347,  -12'd192,  -12'd332,  
12'd548,  12'd135,  -12'd86,  -12'd136,  -12'd104,  -12'd185,  12'd461,  -12'd120,  12'd318,  -12'd125,  12'd185,  12'd101,  12'd538,  12'd203,  -12'd131,  12'd182,  
12'd110,  12'd50,  12'd73,  -12'd154,  12'd290,  -12'd128,  -12'd160,  12'd53,  -12'd245,  -12'd300,  12'd0,  12'd122,  -12'd399,  -12'd5,  -12'd36,  12'd78,  
12'd250,  12'd269,  12'd113,  -12'd21,  12'd68,  -12'd23,  -12'd49,  12'd336,  -12'd386,  -12'd125,  12'd25,  -12'd176,  -12'd125,  -12'd10,  12'd28,  -12'd127,  
12'd171,  12'd396,  -12'd294,  -12'd161,  12'd15,  12'd375,  12'd50,  12'd114,  12'd227,  12'd198,  12'd94,  -12'd295,  12'd374,  -12'd376,  -12'd256,  -12'd416,  
12'd50,  -12'd97,  12'd126,  12'd453,  12'd95,  12'd228,  -12'd196,  12'd321,  -12'd102,  -12'd76,  12'd43,  -12'd200,  -12'd21,  12'd103,  12'd93,  -12'd20,  
12'd657,  12'd395,  -12'd135,  -12'd57,  12'd117,  12'd128,  -12'd218,  -12'd226,  12'd126,  -12'd319,  -12'd145,  12'd46,  12'd482,  -12'd163,  12'd232,  12'd432,  
12'd391,  -12'd282,  -12'd118,  -12'd49,  -12'd262,  -12'd231,  12'd105,  -12'd245,  12'd10,  -12'd246,  -12'd361,  12'd353,  -12'd411,  12'd51,  -12'd177,  12'd15,  
12'd408,  12'd242,  12'd213,  -12'd189,  -12'd141,  12'd54,  12'd166,  -12'd81,  12'd328,  12'd363,  -12'd309,  12'd61,  12'd255,  12'd564,  -12'd127,  12'd45,  
-12'd135,  -12'd16,  -12'd217,  12'd315,  12'd134,  -12'd70,  12'd108,  12'd22,  12'd262,  -12'd21,  12'd210,  12'd55,  -12'd4,  -12'd101,  -12'd281,  12'd72,  
-12'd398,  12'd64,  -12'd403,  -12'd300,  -12'd6,  -12'd267,  -12'd47,  12'd367,  -12'd437,  12'd373,  -12'd128,  -12'd128,  -12'd541,  -12'd137,  -12'd172,  12'd181,  
12'd67,  -12'd285,  -12'd243,  -12'd395,  12'd72,  -12'd223,  -12'd140,  -12'd143,  -12'd288,  -12'd174,  -12'd19,  12'd118,  12'd188,  -12'd61,  -12'd379,  12'd29,  
12'd582,  12'd76,  12'd473,  -12'd205,  -12'd292,  12'd335,  -12'd103,  12'd310,  12'd102,  12'd368,  -12'd2,  12'd323,  12'd40,  12'd577,  12'd255,  12'd293,  
12'd53,  -12'd119,  12'd355,  12'd152,  12'd42,  -12'd394,  -12'd99,  12'd194,  12'd214,  -12'd166,  12'd81,  12'd305,  12'd100,  12'd177,  -12'd119,  -12'd171,  
-12'd273,  12'd66,  -12'd130,  -12'd91,  -12'd68,  -12'd143,  12'd11,  12'd403,  12'd163,  -12'd157,  12'd138,  12'd89,  -12'd60,  12'd262,  12'd12,  -12'd6,  
-12'd193,  -12'd389,  -12'd192,  -12'd148,  12'd310,  -12'd318,  12'd88,  -12'd211,  -12'd469,  12'd40,  -12'd14,  -12'd18,  -12'd245,  -12'd41,  -12'd452,  -12'd167,  
-12'd418,  -12'd565,  12'd154,  -12'd79,  -12'd222,  -12'd92,  -12'd143,  -12'd219,  -12'd220,  -12'd371,  -12'd81,  -12'd185,  12'd86,  -12'd87,  -12'd476,  -12'd126,  

-12'd3,  12'd102,  12'd162,  12'd59,  12'd90,  12'd203,  -12'd306,  12'd245,  -12'd121,  12'd276,  -12'd171,  -12'd180,  12'd67,  12'd76,  12'd91,  12'd76,  
12'd183,  -12'd50,  12'd4,  -12'd24,  12'd298,  12'd232,  -12'd303,  12'd7,  -12'd109,  -12'd151,  -12'd297,  -12'd152,  -12'd122,  12'd179,  12'd133,  12'd76,  
12'd141,  -12'd103,  -12'd137,  12'd97,  -12'd68,  -12'd50,  12'd128,  -12'd156,  -12'd79,  -12'd206,  12'd182,  -12'd409,  -12'd314,  -12'd93,  12'd67,  12'd41,  
-12'd278,  -12'd117,  -12'd41,  -12'd339,  -12'd60,  12'd85,  -12'd76,  -12'd73,  -12'd168,  12'd176,  -12'd239,  -12'd217,  -12'd87,  12'd193,  12'd220,  -12'd312,  
12'd170,  -12'd400,  -12'd195,  -12'd225,  -12'd48,  12'd64,  -12'd203,  -12'd191,  12'd56,  12'd107,  12'd130,  -12'd334,  -12'd289,  -12'd27,  -12'd236,  12'd322,  
-12'd216,  -12'd308,  12'd115,  -12'd96,  -12'd176,  12'd9,  -12'd101,  12'd104,  12'd78,  12'd279,  -12'd106,  12'd151,  12'd83,  -12'd269,  -12'd15,  12'd25,  
12'd70,  -12'd9,  -12'd168,  -12'd311,  -12'd370,  12'd341,  12'd17,  12'd24,  -12'd254,  12'd45,  12'd17,  -12'd170,  -12'd78,  -12'd121,  -12'd234,  12'd89,  
-12'd397,  -12'd252,  12'd43,  -12'd298,  -12'd45,  -12'd107,  -12'd228,  12'd143,  12'd13,  -12'd244,  -12'd100,  -12'd107,  -12'd48,  -12'd135,  12'd350,  -12'd103,  
12'd71,  -12'd75,  -12'd112,  -12'd261,  12'd70,  -12'd187,  -12'd316,  -12'd243,  -12'd162,  -12'd286,  12'd359,  -12'd268,  -12'd315,  -12'd128,  -12'd201,  -12'd71,  
-12'd299,  -12'd35,  12'd151,  -12'd177,  -12'd18,  -12'd116,  -12'd343,  12'd310,  -12'd202,  12'd83,  -12'd40,  -12'd269,  -12'd391,  -12'd82,  -12'd325,  12'd7,  
-12'd266,  -12'd15,  12'd31,  -12'd153,  12'd259,  -12'd83,  -12'd153,  -12'd25,  12'd72,  -12'd276,  12'd30,  12'd13,  -12'd298,  12'd334,  -12'd118,  -12'd60,  
-12'd13,  -12'd369,  -12'd164,  -12'd256,  12'd29,  -12'd64,  12'd86,  -12'd291,  12'd227,  -12'd248,  -12'd156,  12'd334,  -12'd157,  -12'd72,  -12'd18,  12'd114,  
-12'd231,  12'd269,  -12'd5,  -12'd167,  12'd131,  12'd94,  12'd80,  12'd75,  -12'd385,  12'd58,  -12'd104,  -12'd131,  12'd68,  -12'd145,  12'd103,  12'd115,  
-12'd51,  12'd36,  -12'd230,  -12'd341,  12'd246,  -12'd77,  -12'd219,  -12'd114,  -12'd8,  -12'd423,  -12'd235,  -12'd182,  -12'd234,  -12'd267,  -12'd165,  12'd220,  
-12'd144,  12'd204,  -12'd216,  12'd323,  12'd212,  -12'd104,  12'd146,  12'd18,  -12'd200,  -12'd140,  12'd228,  12'd48,  -12'd95,  -12'd116,  -12'd154,  12'd105,  
12'd80,  12'd9,  12'd143,  12'd57,  12'd47,  12'd221,  -12'd124,  -12'd103,  -12'd92,  -12'd384,  -12'd103,  -12'd83,  -12'd355,  -12'd232,  12'd88,  12'd306,  
-12'd150,  -12'd45,  -12'd14,  -12'd265,  12'd158,  -12'd96,  -12'd32,  12'd54,  -12'd89,  -12'd91,  12'd224,  -12'd318,  12'd300,  -12'd308,  -12'd229,  12'd351,  
12'd139,  -12'd32,  -12'd216,  12'd58,  -12'd297,  -12'd196,  -12'd175,  12'd95,  12'd38,  -12'd2,  -12'd347,  -12'd196,  -12'd136,  12'd103,  -12'd236,  -12'd108,  
-12'd224,  -12'd1,  -12'd255,  12'd204,  -12'd127,  -12'd286,  12'd160,  12'd188,  12'd103,  -12'd141,  -12'd47,  -12'd54,  12'd228,  12'd173,  -12'd273,  -12'd208,  
-12'd171,  12'd103,  -12'd148,  -12'd160,  -12'd299,  -12'd85,  12'd150,  -12'd293,  -12'd45,  -12'd107,  -12'd106,  12'd108,  -12'd5,  12'd147,  12'd71,  -12'd339,  
12'd53,  -12'd77,  -12'd165,  -12'd311,  -12'd35,  -12'd118,  12'd315,  12'd29,  12'd373,  12'd59,  -12'd183,  12'd132,  -12'd150,  -12'd106,  -12'd6,  12'd63,  
-12'd3,  12'd107,  -12'd203,  -12'd135,  -12'd127,  12'd223,  12'd43,  12'd227,  12'd92,  12'd68,  12'd152,  12'd107,  12'd32,  -12'd50,  12'd86,  12'd151,  
-12'd71,  -12'd121,  -12'd103,  12'd42,  12'd8,  12'd24,  12'd30,  12'd160,  12'd50,  12'd66,  12'd203,  12'd125,  -12'd345,  -12'd51,  12'd67,  -12'd101,  
12'd153,  -12'd222,  -12'd327,  -12'd418,  -12'd281,  -12'd171,  -12'd117,  -12'd135,  -12'd162,  12'd40,  -12'd80,  -12'd290,  12'd129,  -12'd370,  -12'd187,  -12'd53,  
12'd312,  12'd63,  12'd40,  -12'd83,  12'd76,  -12'd169,  -12'd181,  -12'd62,  -12'd277,  12'd7,  12'd276,  -12'd9,  -12'd194,  -12'd21,  -12'd278,  12'd169,  

12'd177,  12'd74,  -12'd355,  -12'd185,  -12'd547,  -12'd277,  12'd486,  -12'd569,  12'd14,  -12'd279,  -12'd367,  -12'd352,  -12'd238,  12'd216,  -12'd471,  -12'd287,  
12'd236,  -12'd61,  12'd314,  -12'd80,  -12'd71,  -12'd96,  12'd72,  12'd175,  -12'd296,  -12'd267,  -12'd360,  -12'd161,  -12'd320,  12'd360,  12'd56,  -12'd556,  
12'd206,  12'd228,  12'd199,  12'd231,  12'd57,  -12'd318,  12'd138,  12'd164,  12'd88,  12'd67,  12'd281,  12'd72,  12'd106,  -12'd348,  -12'd220,  -12'd510,  
12'd5,  12'd206,  12'd62,  12'd432,  -12'd555,  12'd122,  12'd293,  12'd301,  12'd147,  12'd61,  12'd290,  12'd50,  12'd102,  12'd27,  12'd205,  -12'd324,  
-12'd80,  12'd176,  -12'd13,  12'd511,  -12'd61,  12'd139,  12'd70,  12'd166,  -12'd105,  -12'd96,  12'd155,  -12'd173,  12'd235,  12'd31,  -12'd49,  12'd16,  
-12'd404,  -12'd391,  -12'd277,  -12'd230,  -12'd414,  -12'd437,  12'd111,  -12'd451,  -12'd232,  12'd75,  12'd116,  -12'd266,  -12'd16,  12'd112,  -12'd240,  -12'd364,  
12'd218,  -12'd66,  12'd324,  -12'd213,  -12'd293,  12'd239,  -12'd15,  12'd171,  12'd4,  -12'd74,  -12'd136,  -12'd137,  12'd96,  12'd444,  -12'd38,  -12'd38,  
-12'd224,  -12'd120,  12'd131,  -12'd61,  -12'd13,  12'd157,  12'd142,  12'd447,  12'd376,  12'd244,  12'd180,  -12'd53,  -12'd170,  -12'd543,  12'd77,  -12'd126,  
-12'd155,  12'd17,  12'd89,  12'd463,  12'd251,  -12'd89,  12'd96,  12'd277,  12'd240,  12'd315,  12'd145,  -12'd352,  12'd418,  12'd25,  -12'd159,  12'd193,  
-12'd414,  -12'd47,  -12'd232,  -12'd119,  -12'd4,  -12'd160,  -12'd551,  -12'd139,  -12'd323,  12'd194,  12'd346,  12'd129,  12'd146,  -12'd172,  12'd144,  12'd91,  
-12'd13,  -12'd524,  12'd255,  -12'd115,  -12'd74,  12'd131,  -12'd354,  12'd162,  12'd192,  -12'd239,  -12'd232,  12'd99,  -12'd190,  12'd431,  -12'd72,  -12'd201,  
-12'd21,  -12'd387,  12'd603,  -12'd232,  -12'd286,  12'd68,  12'd112,  12'd0,  -12'd320,  -12'd41,  12'd76,  -12'd1,  12'd24,  12'd2,  12'd114,  12'd189,  
-12'd245,  -12'd80,  12'd5,  -12'd75,  -12'd135,  12'd45,  12'd72,  12'd23,  -12'd327,  12'd169,  -12'd157,  -12'd210,  12'd221,  -12'd110,  12'd123,  -12'd29,  
-12'd508,  -12'd263,  12'd512,  -12'd241,  -12'd43,  -12'd354,  -12'd34,  -12'd33,  -12'd21,  12'd2,  12'd134,  12'd189,  -12'd422,  12'd81,  -12'd1,  -12'd74,  
-12'd668,  12'd439,  12'd87,  -12'd19,  12'd13,  12'd131,  -12'd20,  -12'd8,  12'd16,  -12'd63,  12'd289,  -12'd194,  -12'd709,  -12'd158,  -12'd172,  -12'd300,  
-12'd99,  12'd97,  -12'd316,  -12'd68,  12'd388,  12'd120,  -12'd687,  -12'd202,  -12'd138,  12'd54,  -12'd193,  -12'd246,  -12'd170,  12'd3,  -12'd14,  -12'd251,  
12'd38,  -12'd232,  12'd150,  12'd258,  12'd159,  -12'd122,  -12'd176,  -12'd90,  -12'd647,  -12'd52,  -12'd420,  12'd139,  -12'd84,  12'd133,  12'd29,  12'd81,  
12'd218,  12'd86,  12'd226,  -12'd32,  -12'd173,  12'd47,  12'd327,  -12'd5,  -12'd71,  -12'd227,  -12'd290,  -12'd61,  12'd103,  12'd360,  12'd219,  -12'd33,  
-12'd355,  -12'd194,  12'd409,  12'd259,  -12'd43,  -12'd159,  12'd302,  12'd414,  12'd146,  -12'd214,  -12'd19,  -12'd164,  -12'd138,  -12'd186,  -12'd182,  -12'd87,  
-12'd47,  12'd126,  12'd549,  -12'd433,  -12'd133,  -12'd98,  -12'd197,  12'd149,  -12'd34,  -12'd264,  -12'd90,  -12'd321,  -12'd125,  12'd144,  -12'd274,  -12'd358,  
-12'd458,  12'd54,  -12'd314,  12'd376,  12'd64,  12'd55,  12'd57,  12'd213,  12'd329,  12'd61,  12'd262,  -12'd112,  12'd94,  -12'd513,  12'd28,  -12'd101,  
12'd113,  -12'd117,  12'd19,  12'd230,  12'd219,  -12'd77,  -12'd178,  -12'd195,  12'd330,  12'd1,  12'd423,  -12'd54,  12'd103,  -12'd489,  -12'd31,  -12'd36,  
12'd244,  12'd247,  12'd269,  -12'd6,  12'd188,  12'd45,  -12'd170,  12'd24,  -12'd146,  12'd328,  12'd26,  12'd68,  -12'd341,  12'd356,  12'd108,  -12'd78,  
-12'd399,  12'd9,  12'd56,  12'd325,  -12'd272,  -12'd178,  12'd319,  -12'd60,  -12'd190,  -12'd289,  12'd175,  -12'd179,  -12'd125,  -12'd320,  12'd28,  -12'd119,  
-12'd243,  -12'd465,  -12'd418,  -12'd190,  -12'd430,  -12'd659,  12'd205,  -12'd289,  12'd176,  -12'd45,  -12'd325,  -12'd79,  -12'd162,  12'd191,  -12'd112,  -12'd403,  

12'd19,  12'd115,  12'd317,  12'd234,  -12'd167,  -12'd402,  12'd157,  -12'd42,  -12'd127,  -12'd17,  12'd264,  -12'd296,  -12'd153,  -12'd2,  -12'd314,  -12'd64,  
12'd176,  -12'd63,  -12'd50,  -12'd65,  -12'd393,  12'd235,  12'd91,  -12'd179,  -12'd111,  -12'd310,  12'd139,  -12'd203,  -12'd71,  -12'd309,  -12'd332,  12'd143,  
-12'd97,  12'd142,  12'd49,  12'd155,  -12'd314,  -12'd218,  -12'd22,  -12'd213,  12'd11,  -12'd175,  12'd113,  12'd171,  -12'd55,  12'd124,  12'd78,  12'd5,  
-12'd143,  12'd202,  -12'd260,  12'd14,  12'd230,  -12'd441,  12'd104,  -12'd16,  -12'd169,  -12'd282,  12'd281,  12'd50,  12'd0,  -12'd115,  12'd155,  12'd26,  
12'd151,  12'd173,  -12'd195,  -12'd23,  12'd265,  -12'd77,  -12'd139,  -12'd52,  12'd74,  12'd119,  12'd304,  -12'd230,  -12'd12,  12'd214,  -12'd223,  12'd231,  
-12'd292,  -12'd185,  12'd97,  -12'd28,  -12'd211,  -12'd159,  12'd128,  -12'd53,  -12'd68,  12'd185,  12'd149,  -12'd190,  -12'd185,  12'd119,  -12'd128,  12'd8,  
12'd138,  -12'd128,  -12'd12,  -12'd227,  -12'd217,  -12'd28,  -12'd183,  -12'd179,  -12'd93,  -12'd27,  12'd288,  -12'd134,  -12'd212,  12'd112,  12'd34,  -12'd155,  
-12'd80,  12'd83,  -12'd156,  -12'd243,  12'd197,  -12'd84,  -12'd144,  -12'd242,  -12'd36,  12'd12,  -12'd63,  12'd151,  -12'd195,  12'd349,  -12'd404,  -12'd378,  
-12'd323,  12'd129,  -12'd287,  12'd88,  -12'd62,  -12'd172,  -12'd188,  12'd161,  -12'd161,  -12'd299,  -12'd431,  -12'd31,  -12'd7,  12'd56,  -12'd6,  12'd48,  
12'd56,  12'd276,  -12'd123,  12'd156,  -12'd261,  -12'd86,  -12'd2,  -12'd271,  12'd290,  -12'd76,  12'd37,  -12'd316,  -12'd36,  12'd76,  12'd237,  -12'd160,  
-12'd292,  12'd78,  12'd145,  -12'd323,  12'd36,  -12'd32,  -12'd312,  12'd163,  -12'd63,  12'd82,  -12'd184,  -12'd141,  12'd54,  -12'd295,  -12'd166,  -12'd4,  
-12'd231,  -12'd403,  -12'd5,  -12'd84,  -12'd408,  -12'd312,  -12'd145,  -12'd347,  -12'd155,  -12'd139,  -12'd22,  12'd196,  12'd40,  -12'd34,  -12'd77,  12'd132,  
-12'd112,  -12'd109,  12'd221,  -12'd197,  -12'd323,  -12'd289,  12'd96,  -12'd31,  -12'd11,  -12'd164,  -12'd244,  -12'd402,  -12'd36,  -12'd42,  -12'd146,  -12'd77,  
12'd20,  12'd166,  -12'd248,  12'd290,  -12'd231,  -12'd60,  -12'd259,  -12'd145,  12'd112,  -12'd7,  -12'd97,  -12'd154,  12'd105,  12'd121,  -12'd27,  12'd172,  
-12'd109,  12'd104,  -12'd15,  -12'd112,  12'd4,  12'd29,  -12'd114,  12'd117,  -12'd244,  -12'd88,  -12'd364,  -12'd363,  12'd76,  12'd255,  12'd33,  12'd107,  
-12'd105,  12'd20,  -12'd54,  12'd267,  12'd215,  -12'd18,  -12'd89,  -12'd184,  12'd83,  -12'd163,  12'd250,  12'd260,  -12'd57,  -12'd103,  -12'd250,  12'd168,  
12'd84,  -12'd9,  -12'd227,  -12'd1,  12'd13,  -12'd322,  -12'd18,  12'd104,  12'd105,  -12'd79,  -12'd235,  -12'd159,  -12'd238,  -12'd56,  -12'd161,  12'd148,  
12'd142,  -12'd10,  -12'd228,  12'd213,  12'd52,  12'd78,  12'd45,  12'd21,  -12'd90,  12'd297,  12'd360,  -12'd359,  -12'd56,  -12'd24,  -12'd235,  12'd15,  
-12'd101,  -12'd82,  -12'd89,  -12'd241,  -12'd276,  -12'd202,  -12'd228,  -12'd40,  -12'd301,  12'd59,  12'd174,  -12'd408,  12'd204,  -12'd412,  12'd55,  -12'd211,  
12'd371,  -12'd97,  12'd119,  -12'd123,  12'd109,  -12'd325,  -12'd291,  -12'd352,  -12'd123,  12'd95,  12'd190,  12'd279,  -12'd216,  12'd8,  -12'd151,  12'd32,  
-12'd41,  12'd38,  12'd99,  -12'd42,  12'd27,  12'd331,  -12'd70,  12'd9,  -12'd70,  -12'd314,  12'd157,  -12'd119,  12'd40,  12'd142,  12'd51,  -12'd92,  
-12'd340,  -12'd147,  -12'd146,  -12'd75,  12'd116,  12'd50,  -12'd2,  12'd51,  -12'd253,  -12'd235,  12'd143,  12'd89,  12'd280,  12'd165,  -12'd397,  12'd126,  
-12'd117,  -12'd47,  12'd178,  -12'd423,  -12'd283,  -12'd424,  -12'd20,  12'd239,  -12'd168,  -12'd231,  12'd53,  12'd66,  -12'd161,  -12'd81,  12'd315,  12'd34,  
-12'd19,  -12'd246,  12'd267,  -12'd53,  -12'd304,  -12'd171,  12'd67,  12'd46,  -12'd1,  -12'd50,  -12'd294,  -12'd150,  12'd248,  12'd55,  12'd41,  12'd127,  
-12'd87,  -12'd257,  12'd84,  12'd178,  -12'd7,  12'd28,  -12'd12,  12'd35,  -12'd66,  -12'd109,  -12'd139,  12'd70,  12'd144,  -12'd192,  12'd129,  12'd102,  

-12'd103,  -12'd393,  12'd35,  12'd39,  -12'd32,  -12'd161,  12'd285,  12'd391,  12'd206,  12'd78,  12'd148,  -12'd423,  12'd170,  -12'd175,  12'd197,  12'd77,  
12'd256,  12'd80,  -12'd2,  -12'd304,  12'd286,  -12'd22,  -12'd44,  12'd411,  -12'd75,  12'd298,  12'd251,  -12'd28,  12'd425,  -12'd278,  12'd199,  -12'd374,  
12'd3,  -12'd305,  12'd62,  12'd228,  -12'd268,  12'd140,  12'd1,  -12'd70,  12'd0,  12'd10,  -12'd66,  12'd153,  12'd332,  -12'd202,  12'd11,  -12'd45,  
12'd460,  -12'd12,  12'd298,  -12'd36,  -12'd188,  -12'd278,  12'd116,  12'd66,  12'd330,  -12'd296,  12'd14,  -12'd170,  12'd490,  -12'd237,  12'd404,  -12'd37,  
-12'd134,  -12'd227,  12'd130,  -12'd303,  -12'd86,  -12'd209,  -12'd265,  12'd324,  12'd27,  -12'd50,  12'd215,  12'd206,  12'd205,  -12'd207,  -12'd184,  12'd3,  
-12'd29,  12'd206,  12'd170,  12'd279,  12'd373,  -12'd177,  -12'd427,  -12'd157,  -12'd56,  -12'd38,  -12'd59,  12'd36,  -12'd47,  -12'd17,  -12'd353,  -12'd52,  
-12'd358,  12'd438,  12'd32,  -12'd148,  -12'd163,  12'd258,  -12'd254,  -12'd252,  12'd275,  -12'd28,  -12'd77,  -12'd86,  12'd3,  -12'd3,  -12'd240,  -12'd203,  
-12'd366,  12'd411,  -12'd102,  12'd116,  12'd230,  12'd184,  12'd39,  -12'd0,  -12'd117,  12'd100,  12'd240,  -12'd100,  12'd192,  12'd94,  12'd132,  12'd390,  
-12'd171,  12'd364,  -12'd24,  12'd13,  12'd128,  -12'd217,  -12'd293,  -12'd26,  12'd85,  -12'd198,  12'd144,  -12'd33,  12'd227,  12'd72,  12'd154,  12'd84,  
-12'd193,  12'd111,  12'd85,  12'd167,  -12'd249,  12'd129,  -12'd351,  -12'd241,  -12'd57,  12'd165,  -12'd225,  12'd536,  12'd267,  -12'd120,  12'd151,  12'd345,  
-12'd84,  12'd63,  12'd7,  -12'd252,  -12'd3,  -12'd41,  -12'd272,  12'd20,  12'd230,  -12'd252,  12'd565,  12'd224,  12'd82,  12'd12,  12'd194,  -12'd264,  
12'd271,  12'd218,  12'd445,  -12'd316,  -12'd124,  -12'd199,  -12'd30,  -12'd326,  12'd198,  12'd37,  12'd35,  -12'd25,  -12'd264,  -12'd17,  -12'd271,  12'd215,  
12'd95,  12'd59,  -12'd134,  12'd2,  -12'd55,  -12'd113,  12'd50,  -12'd63,  -12'd169,  -12'd94,  12'd8,  -12'd275,  12'd55,  12'd139,  12'd45,  12'd4,  
-12'd225,  12'd169,  -12'd211,  -12'd203,  12'd477,  12'd234,  12'd28,  -12'd272,  -12'd193,  12'd84,  12'd75,  12'd191,  12'd222,  -12'd15,  -12'd22,  12'd31,  
12'd35,  12'd122,  12'd694,  12'd128,  12'd410,  -12'd427,  12'd111,  12'd24,  12'd160,  12'd356,  12'd209,  12'd294,  -12'd190,  12'd8,  12'd26,  12'd341,  
12'd323,  12'd103,  12'd101,  -12'd239,  -12'd69,  -12'd346,  12'd174,  12'd11,  -12'd70,  -12'd233,  12'd227,  -12'd99,  -12'd286,  12'd41,  12'd42,  12'd0,  
12'd307,  12'd44,  12'd21,  12'd24,  12'd101,  -12'd224,  12'd234,  -12'd131,  12'd101,  12'd151,  -12'd157,  12'd117,  12'd155,  12'd293,  -12'd182,  -12'd74,  
-12'd87,  -12'd71,  12'd132,  -12'd327,  -12'd127,  12'd220,  12'd175,  12'd67,  12'd159,  -12'd350,  -12'd44,  12'd376,  12'd24,  -12'd172,  -12'd148,  -12'd221,  
-12'd50,  -12'd237,  12'd2,  -12'd60,  -12'd228,  12'd186,  12'd234,  -12'd106,  -12'd105,  -12'd113,  -12'd141,  12'd125,  12'd103,  12'd95,  -12'd413,  12'd14,  
-12'd130,  12'd25,  12'd372,  12'd142,  -12'd386,  12'd85,  12'd245,  12'd207,  12'd144,  -12'd185,  -12'd95,  -12'd111,  12'd291,  -12'd113,  12'd200,  -12'd269,  
-12'd107,  -12'd20,  12'd90,  12'd134,  -12'd153,  -12'd76,  -12'd24,  12'd259,  -12'd87,  -12'd34,  -12'd262,  -12'd303,  12'd101,  12'd314,  -12'd106,  12'd277,  
12'd70,  -12'd7,  12'd191,  12'd167,  -12'd212,  12'd174,  -12'd302,  12'd314,  -12'd268,  12'd290,  12'd59,  12'd200,  12'd110,  12'd124,  12'd454,  -12'd49,  
12'd294,  12'd79,  -12'd131,  12'd29,  12'd79,  12'd163,  -12'd155,  -12'd249,  12'd190,  -12'd151,  12'd290,  12'd105,  12'd60,  -12'd49,  -12'd258,  -12'd98,  
12'd59,  -12'd107,  12'd172,  -12'd358,  12'd73,  -12'd119,  12'd279,  -12'd170,  -12'd218,  12'd27,  -12'd15,  12'd141,  -12'd132,  12'd115,  -12'd48,  12'd132,  
12'd193,  12'd105,  12'd402,  -12'd293,  -12'd298,  -12'd47,  12'd1,  -12'd54,  12'd43,  -12'd50,  -12'd250,  -12'd140,  -12'd434,  12'd330,  -12'd204,  -12'd144,  

12'd51,  12'd259,  12'd132,  -12'd61,  12'd95,  12'd68,  12'd269,  12'd131,  -12'd88,  -12'd12,  12'd101,  -12'd1,  12'd157,  12'd166,  12'd352,  -12'd3,  
12'd524,  12'd108,  12'd418,  -12'd113,  -12'd242,  12'd118,  12'd372,  -12'd189,  -12'd7,  -12'd308,  12'd251,  12'd184,  -12'd20,  12'd397,  -12'd117,  12'd286,  
12'd144,  -12'd107,  12'd347,  -12'd198,  -12'd287,  -12'd217,  12'd517,  -12'd369,  -12'd426,  -12'd214,  12'd154,  -12'd374,  12'd65,  12'd80,  -12'd361,  -12'd178,  
-12'd194,  -12'd11,  -12'd672,  -12'd513,  -12'd41,  -12'd339,  12'd473,  -12'd366,  -12'd262,  -12'd563,  12'd443,  -12'd11,  -12'd80,  12'd293,  -12'd209,  -12'd43,  
-12'd244,  12'd72,  -12'd550,  -12'd296,  -12'd339,  -12'd220,  -12'd568,  -12'd549,  -12'd493,  -12'd139,  -12'd30,  -12'd352,  -12'd520,  -12'd80,  -12'd275,  12'd233,  
12'd427,  -12'd30,  12'd144,  -12'd3,  -12'd204,  -12'd238,  12'd14,  12'd16,  12'd361,  -12'd300,  12'd341,  12'd326,  12'd498,  12'd26,  12'd222,  12'd64,  
-12'd15,  12'd284,  -12'd110,  -12'd301,  12'd207,  -12'd276,  12'd211,  12'd4,  -12'd260,  12'd305,  12'd238,  -12'd151,  -12'd35,  12'd136,  12'd39,  12'd36,  
-12'd78,  -12'd399,  12'd144,  -12'd152,  -12'd154,  -12'd732,  -12'd49,  -12'd288,  12'd87,  -12'd18,  12'd55,  12'd177,  -12'd89,  -12'd261,  -12'd354,  -12'd354,  
12'd87,  12'd84,  -12'd283,  -12'd46,  -12'd282,  12'd63,  -12'd157,  -12'd547,  12'd413,  12'd356,  -12'd194,  -12'd237,  -12'd151,  -12'd180,  -12'd309,  -12'd341,  
12'd418,  -12'd452,  -12'd6,  12'd251,  12'd313,  -12'd106,  -12'd3,  -12'd451,  12'd119,  12'd343,  -12'd337,  12'd442,  12'd45,  12'd17,  -12'd198,  12'd39,  
-12'd191,  12'd13,  12'd336,  12'd69,  -12'd225,  -12'd250,  12'd187,  -12'd55,  -12'd115,  12'd17,  -12'd2,  -12'd149,  -12'd324,  12'd5,  -12'd267,  12'd164,  
-12'd306,  12'd358,  12'd438,  -12'd304,  -12'd144,  -12'd189,  12'd67,  -12'd74,  12'd112,  -12'd173,  -12'd237,  -12'd362,  -12'd353,  12'd313,  12'd62,  -12'd544,  
12'd237,  -12'd599,  12'd211,  12'd46,  -12'd333,  -12'd228,  -12'd344,  -12'd240,  -12'd265,  12'd96,  -12'd244,  -12'd26,  -12'd608,  -12'd16,  -12'd148,  12'd90,  
12'd412,  -12'd141,  -12'd528,  12'd134,  12'd18,  12'd244,  -12'd244,  -12'd51,  12'd444,  12'd76,  12'd456,  12'd211,  12'd183,  -12'd9,  -12'd63,  12'd278,  
12'd280,  12'd159,  12'd78,  12'd127,  12'd350,  12'd326,  12'd236,  -12'd55,  12'd258,  12'd253,  12'd553,  12'd289,  12'd187,  -12'd51,  12'd239,  12'd171,  
-12'd207,  12'd108,  -12'd293,  -12'd2,  12'd252,  -12'd154,  12'd90,  12'd148,  12'd173,  -12'd420,  -12'd183,  -12'd206,  12'd212,  -12'd93,  12'd113,  12'd132,  
12'd29,  -12'd190,  12'd158,  12'd132,  -12'd154,  12'd277,  -12'd128,  12'd164,  -12'd158,  -12'd52,  12'd211,  -12'd63,  12'd32,  12'd324,  12'd13,  -12'd190,  
12'd137,  -12'd381,  12'd302,  12'd267,  -12'd80,  -12'd90,  -12'd109,  12'd259,  -12'd532,  12'd90,  12'd232,  -12'd42,  12'd402,  -12'd140,  12'd196,  -12'd508,  
-12'd18,  -12'd140,  -12'd252,  12'd384,  12'd366,  -12'd7,  12'd275,  12'd235,  -12'd430,  -12'd150,  12'd307,  12'd204,  12'd179,  -12'd209,  12'd369,  -12'd13,  
-12'd55,  12'd34,  -12'd135,  12'd205,  -12'd127,  12'd49,  12'd176,  12'd438,  -12'd186,  12'd309,  12'd191,  12'd74,  12'd452,  -12'd68,  12'd56,  12'd194,  
12'd49,  -12'd49,  12'd37,  12'd12,  12'd233,  -12'd164,  -12'd468,  12'd131,  12'd70,  12'd49,  12'd16,  -12'd515,  12'd122,  -12'd25,  -12'd337,  -12'd140,  
-12'd432,  12'd203,  -12'd146,  12'd183,  -12'd132,  -12'd28,  -12'd692,  12'd127,  12'd375,  12'd83,  12'd158,  -12'd591,  12'd255,  12'd229,  -12'd262,  12'd120,  
12'd9,  -12'd177,  -12'd603,  12'd47,  -12'd229,  12'd243,  -12'd111,  12'd71,  -12'd511,  -12'd113,  12'd327,  12'd5,  12'd300,  -12'd902,  -12'd273,  -12'd210,  
-12'd419,  -12'd381,  -12'd1005,  12'd32,  12'd201,  -12'd96,  -12'd116,  -12'd27,  12'd145,  -12'd468,  12'd247,  12'd7,  12'd34,  -12'd42,  -12'd398,  12'd1,  
12'd38,  -12'd416,  -12'd338,  -12'd364,  12'd87,  -12'd528,  -12'd344,  12'd234,  -12'd74,  12'd508,  12'd9,  -12'd318,  -12'd301,  -12'd236,  -12'd227,  12'd184,  

-12'd169,  -12'd146,  12'd329,  12'd227,  -12'd62,  -12'd129,  -12'd295,  12'd91,  12'd69,  -12'd98,  -12'd151,  -12'd121,  -12'd164,  -12'd158,  12'd162,  -12'd86,  
12'd379,  -12'd231,  12'd157,  12'd403,  12'd112,  12'd429,  -12'd82,  12'd119,  -12'd222,  -12'd235,  -12'd298,  12'd29,  12'd356,  12'd146,  12'd252,  -12'd544,  
-12'd165,  12'd99,  -12'd92,  -12'd136,  -12'd112,  12'd459,  -12'd160,  12'd303,  12'd596,  12'd295,  -12'd16,  -12'd305,  12'd271,  -12'd256,  12'd415,  -12'd288,  
-12'd39,  -12'd116,  -12'd238,  12'd56,  -12'd210,  -12'd209,  -12'd503,  -12'd15,  -12'd431,  12'd187,  -12'd241,  -12'd324,  12'd1,  -12'd343,  12'd121,  12'd393,  
-12'd30,  -12'd199,  12'd177,  12'd42,  12'd140,  -12'd47,  12'd147,  12'd315,  -12'd23,  12'd141,  -12'd21,  12'd125,  12'd13,  -12'd203,  -12'd54,  -12'd327,  
12'd246,  -12'd40,  12'd59,  -12'd191,  -12'd298,  12'd92,  12'd40,  -12'd128,  -12'd108,  12'd46,  -12'd32,  12'd199,  -12'd110,  12'd322,  12'd244,  -12'd199,  
12'd159,  -12'd266,  12'd685,  12'd139,  -12'd38,  12'd364,  -12'd184,  12'd64,  12'd251,  -12'd384,  -12'd335,  -12'd329,  -12'd63,  12'd18,  -12'd339,  -12'd208,  
-12'd207,  12'd505,  -12'd354,  -12'd211,  12'd130,  12'd580,  -12'd96,  12'd390,  12'd435,  -12'd150,  -12'd5,  12'd52,  12'd156,  12'd171,  12'd21,  12'd137,  
12'd125,  12'd162,  -12'd98,  12'd76,  12'd71,  12'd136,  -12'd299,  12'd273,  -12'd289,  -12'd27,  -12'd127,  -12'd301,  12'd220,  12'd124,  12'd360,  -12'd179,  
-12'd43,  -12'd219,  12'd36,  12'd76,  12'd325,  12'd66,  12'd12,  12'd104,  -12'd227,  12'd185,  12'd361,  12'd578,  12'd57,  -12'd294,  12'd51,  12'd244,  
12'd194,  -12'd146,  12'd359,  12'd236,  12'd57,  12'd363,  -12'd24,  12'd67,  -12'd114,  -12'd86,  -12'd17,  12'd185,  -12'd279,  12'd58,  -12'd222,  -12'd227,  
12'd189,  12'd495,  -12'd11,  -12'd122,  12'd144,  12'd230,  12'd261,  -12'd220,  -12'd2,  -12'd309,  12'd45,  12'd81,  12'd260,  -12'd217,  -12'd257,  -12'd66,  
12'd134,  12'd386,  -12'd375,  12'd58,  12'd320,  -12'd25,  12'd247,  -12'd315,  -12'd217,  -12'd70,  -12'd335,  -12'd503,  -12'd269,  12'd199,  12'd49,  -12'd273,  
12'd208,  12'd448,  -12'd223,  -12'd474,  12'd233,  12'd3,  -12'd188,  12'd14,  -12'd101,  -12'd224,  -12'd209,  12'd55,  -12'd53,  12'd138,  12'd376,  12'd135,  
12'd105,  12'd317,  12'd66,  -12'd39,  12'd287,  -12'd88,  -12'd17,  -12'd88,  -12'd184,  -12'd848,  12'd193,  -12'd176,  12'd2,  -12'd240,  12'd136,  12'd14,  
12'd192,  -12'd145,  12'd128,  12'd310,  12'd36,  -12'd97,  12'd50,  12'd288,  -12'd242,  -12'd140,  -12'd276,  -12'd32,  -12'd254,  -12'd105,  12'd164,  -12'd63,  
12'd9,  -12'd105,  -12'd93,  -12'd286,  -12'd86,  -12'd125,  12'd586,  12'd296,  -12'd49,  -12'd416,  -12'd211,  -12'd117,  -12'd423,  12'd47,  12'd247,  -12'd404,  
12'd251,  12'd157,  12'd211,  12'd122,  -12'd71,  -12'd156,  -12'd81,  -12'd59,  12'd221,  12'd25,  -12'd12,  -12'd39,  -12'd222,  12'd370,  -12'd32,  -12'd309,  
12'd271,  12'd270,  12'd95,  -12'd101,  12'd12,  12'd246,  12'd176,  -12'd52,  12'd5,  12'd131,  12'd108,  12'd267,  12'd135,  12'd358,  -12'd338,  -12'd139,  
12'd206,  12'd198,  12'd267,  -12'd165,  12'd75,  12'd262,  12'd258,  12'd213,  -12'd79,  -12'd109,  12'd57,  12'd111,  -12'd38,  -12'd43,  -12'd504,  12'd128,  
-12'd259,  12'd265,  12'd62,  12'd0,  -12'd351,  12'd144,  -12'd93,  12'd284,  12'd55,  -12'd58,  -12'd71,  12'd284,  -12'd208,  -12'd183,  -12'd213,  12'd49,  
12'd82,  -12'd79,  -12'd189,  -12'd69,  12'd34,  12'd226,  12'd65,  12'd34,  12'd66,  12'd106,  12'd3,  12'd109,  12'd204,  -12'd150,  12'd55,  -12'd69,  
-12'd149,  -12'd371,  -12'd177,  -12'd105,  12'd99,  12'd57,  -12'd142,  -12'd51,  12'd119,  12'd45,  -12'd130,  12'd217,  -12'd25,  -12'd151,  -12'd322,  12'd54,  
12'd619,  -12'd370,  12'd434,  -12'd110,  12'd219,  12'd8,  -12'd185,  12'd129,  12'd176,  12'd136,  12'd234,  12'd290,  12'd107,  -12'd113,  -12'd590,  -12'd234,  
12'd502,  12'd243,  -12'd108,  -12'd483,  -12'd109,  -12'd344,  -12'd247,  12'd46,  -12'd270,  -12'd409,  -12'd438,  -12'd220,  12'd63,  -12'd165,  -12'd559,  12'd128,  

12'd375,  12'd153,  -12'd297,  -12'd12,  -12'd112,  -12'd168,  12'd227,  -12'd170,  12'd295,  -12'd155,  -12'd177,  12'd82,  -12'd512,  -12'd148,  12'd136,  -12'd338,  
12'd261,  12'd150,  12'd47,  -12'd175,  -12'd215,  12'd3,  -12'd85,  12'd225,  -12'd125,  12'd313,  -12'd120,  -12'd170,  -12'd56,  -12'd57,  12'd68,  -12'd88,  
12'd191,  -12'd151,  -12'd90,  12'd22,  12'd7,  12'd56,  -12'd385,  -12'd264,  12'd1,  12'd425,  -12'd34,  12'd21,  -12'd283,  -12'd103,  12'd101,  12'd346,  
-12'd114,  -12'd227,  12'd142,  12'd173,  -12'd142,  -12'd226,  -12'd96,  -12'd164,  12'd141,  12'd75,  12'd257,  -12'd428,  12'd274,  -12'd315,  -12'd61,  12'd24,  
12'd303,  -12'd196,  12'd54,  -12'd14,  12'd398,  -12'd137,  -12'd162,  12'd203,  -12'd218,  -12'd163,  12'd118,  12'd94,  -12'd146,  12'd42,  -12'd9,  12'd574,  
12'd59,  -12'd72,  12'd269,  -12'd81,  12'd323,  12'd157,  -12'd254,  -12'd20,  12'd211,  12'd413,  -12'd234,  -12'd20,  -12'd111,  -12'd184,  12'd490,  12'd55,  
-12'd152,  12'd247,  12'd159,  12'd18,  12'd111,  -12'd124,  -12'd70,  12'd415,  12'd53,  12'd186,  -12'd414,  -12'd236,  12'd106,  12'd170,  12'd390,  12'd524,  
-12'd106,  -12'd6,  12'd57,  12'd278,  -12'd366,  -12'd38,  -12'd178,  12'd134,  12'd71,  -12'd235,  12'd87,  -12'd14,  12'd227,  -12'd296,  -12'd168,  12'd28,  
-12'd249,  -12'd177,  -12'd248,  -12'd13,  -12'd206,  -12'd82,  12'd48,  12'd61,  -12'd72,  12'd61,  -12'd159,  12'd280,  -12'd150,  -12'd489,  -12'd177,  12'd136,  
-12'd8,  12'd378,  -12'd220,  -12'd126,  -12'd0,  12'd188,  -12'd16,  12'd391,  -12'd145,  12'd180,  -12'd154,  12'd167,  12'd454,  12'd22,  -12'd275,  12'd4,  
-12'd133,  -12'd184,  -12'd213,  12'd423,  12'd463,  12'd89,  -12'd928,  12'd317,  -12'd1,  12'd455,  12'd16,  12'd487,  -12'd97,  -12'd147,  -12'd31,  12'd23,  
-12'd105,  12'd617,  12'd237,  12'd61,  -12'd14,  12'd261,  -12'd203,  12'd50,  -12'd74,  12'd391,  12'd441,  12'd259,  -12'd6,  12'd56,  -12'd34,  12'd287,  
12'd109,  12'd15,  -12'd1,  12'd212,  -12'd187,  12'd2,  -12'd317,  -12'd144,  -12'd46,  12'd78,  12'd260,  12'd353,  12'd6,  -12'd264,  -12'd73,  12'd92,  
-12'd293,  -12'd221,  12'd16,  -12'd211,  12'd327,  -12'd408,  12'd192,  12'd98,  -12'd145,  -12'd28,  12'd186,  12'd89,  12'd236,  12'd187,  -12'd25,  12'd384,  
12'd391,  -12'd138,  -12'd353,  -12'd40,  12'd70,  12'd4,  -12'd137,  -12'd355,  -12'd154,  -12'd5,  -12'd34,  -12'd147,  12'd130,  -12'd88,  -12'd107,  12'd201,  
-12'd35,  -12'd324,  -12'd74,  12'd206,  12'd686,  -12'd25,  -12'd351,  12'd125,  12'd146,  12'd234,  -12'd110,  12'd418,  -12'd87,  12'd211,  12'd245,  12'd35,  
12'd246,  12'd135,  -12'd106,  12'd175,  12'd340,  -12'd8,  12'd67,  -12'd426,  12'd430,  12'd490,  -12'd186,  12'd234,  12'd356,  -12'd24,  -12'd66,  12'd143,  
-12'd108,  12'd358,  12'd35,  -12'd132,  12'd83,  -12'd411,  12'd172,  -12'd68,  12'd362,  -12'd168,  -12'd184,  12'd128,  -12'd312,  12'd186,  -12'd161,  -12'd278,  
12'd109,  -12'd41,  12'd36,  -12'd368,  12'd5,  -12'd5,  -12'd284,  -12'd151,  -12'd45,  -12'd86,  -12'd536,  12'd61,  12'd90,  12'd43,  -12'd158,  -12'd393,  
-12'd175,  -12'd39,  12'd439,  -12'd11,  -12'd77,  12'd67,  12'd70,  -12'd84,  12'd101,  12'd37,  -12'd404,  12'd213,  -12'd164,  12'd11,  12'd196,  -12'd399,  
12'd125,  12'd84,  -12'd6,  -12'd39,  12'd67,  12'd385,  12'd296,  12'd493,  12'd168,  -12'd25,  -12'd26,  12'd315,  12'd56,  12'd62,  12'd16,  12'd237,  
-12'd36,  -12'd58,  -12'd273,  12'd138,  -12'd15,  -12'd37,  -12'd500,  12'd311,  -12'd302,  -12'd4,  -12'd51,  -12'd262,  12'd150,  12'd175,  12'd261,  -12'd80,  
12'd216,  -12'd388,  -12'd153,  -12'd96,  -12'd288,  -12'd194,  12'd153,  -12'd82,  12'd57,  12'd393,  12'd28,  12'd464,  12'd108,  -12'd14,  12'd140,  -12'd185,  
12'd46,  -12'd123,  -12'd98,  12'd292,  -12'd176,  12'd359,  -12'd314,  -12'd329,  12'd130,  -12'd14,  12'd279,  12'd314,  -12'd0,  12'd150,  12'd52,  -12'd91,  
12'd394,  -12'd132,  12'd673,  12'd325,  -12'd157,  12'd498,  -12'd42,  12'd144,  12'd399,  -12'd119,  -12'd57,  12'd133,  -12'd59,  12'd3,  12'd413,  -12'd241,  

-12'd130,  12'd183,  -12'd125,  -12'd174,  -12'd51,  12'd96,  12'd97,  12'd297,  12'd235,  -12'd34,  12'd14,  -12'd65,  12'd552,  12'd199,  12'd47,  -12'd87,  
12'd225,  12'd294,  12'd456,  -12'd17,  12'd32,  12'd117,  12'd124,  12'd53,  12'd121,  12'd10,  12'd130,  -12'd307,  12'd175,  12'd88,  12'd127,  12'd215,  
-12'd157,  -12'd181,  12'd103,  12'd160,  -12'd32,  12'd36,  12'd157,  12'd222,  12'd65,  12'd17,  -12'd76,  12'd92,  12'd130,  -12'd103,  -12'd143,  12'd241,  
12'd192,  12'd46,  12'd316,  12'd121,  -12'd261,  12'd149,  -12'd231,  -12'd22,  -12'd120,  -12'd84,  -12'd179,  12'd117,  12'd244,  -12'd175,  -12'd39,  12'd30,  
12'd105,  12'd197,  12'd70,  -12'd98,  -12'd139,  -12'd19,  12'd61,  -12'd4,  -12'd79,  -12'd211,  -12'd200,  12'd250,  -12'd106,  -12'd167,  12'd138,  -12'd313,  
-12'd237,  12'd97,  -12'd168,  12'd137,  12'd19,  12'd74,  -12'd189,  -12'd360,  -12'd89,  -12'd373,  12'd256,  12'd166,  12'd3,  12'd314,  -12'd0,  12'd232,  
-12'd108,  12'd4,  12'd445,  -12'd204,  -12'd185,  12'd345,  12'd255,  -12'd468,  -12'd4,  -12'd146,  12'd366,  12'd28,  12'd39,  12'd173,  -12'd308,  12'd84,  
12'd11,  12'd563,  -12'd282,  12'd209,  12'd135,  12'd383,  12'd555,  -12'd236,  12'd43,  12'd84,  12'd33,  -12'd25,  -12'd90,  12'd216,  -12'd65,  12'd393,  
12'd1,  12'd344,  12'd53,  -12'd274,  12'd445,  -12'd100,  -12'd150,  12'd131,  -12'd219,  12'd229,  -12'd28,  12'd27,  12'd312,  -12'd169,  12'd106,  12'd49,  
12'd597,  12'd124,  -12'd159,  -12'd391,  -12'd151,  -12'd212,  -12'd38,  -12'd200,  12'd324,  12'd465,  12'd66,  12'd249,  -12'd83,  -12'd260,  12'd114,  12'd15,  
-12'd87,  -12'd178,  -12'd82,  -12'd194,  -12'd390,  -12'd222,  12'd196,  12'd229,  -12'd151,  -12'd40,  12'd143,  12'd170,  12'd186,  -12'd120,  12'd43,  -12'd78,  
12'd303,  12'd112,  12'd19,  -12'd185,  12'd16,  -12'd268,  12'd186,  -12'd172,  -12'd274,  -12'd281,  -12'd112,  -12'd123,  12'd12,  12'd36,  12'd64,  -12'd18,  
-12'd8,  12'd593,  12'd164,  -12'd346,  12'd149,  -12'd321,  12'd287,  -12'd20,  -12'd68,  12'd187,  -12'd393,  -12'd101,  -12'd625,  12'd609,  -12'd3,  12'd256,  
-12'd148,  12'd295,  12'd245,  -12'd92,  12'd26,  -12'd98,  12'd92,  12'd208,  12'd19,  -12'd283,  12'd35,  12'd29,  -12'd552,  12'd238,  12'd69,  -12'd367,  
12'd41,  12'd43,  12'd253,  -12'd437,  -12'd393,  -12'd21,  12'd256,  -12'd12,  -12'd87,  -12'd253,  -12'd225,  -12'd108,  -12'd231,  -12'd231,  12'd515,  -12'd371,  
12'd568,  12'd44,  12'd62,  -12'd590,  -12'd258,  -12'd193,  12'd19,  -12'd362,  -12'd237,  12'd13,  -12'd392,  12'd270,  -12'd665,  12'd142,  -12'd202,  12'd166,  
-12'd126,  12'd260,  12'd217,  -12'd275,  -12'd368,  -12'd110,  12'd274,  -12'd46,  12'd639,  12'd246,  -12'd41,  12'd170,  -12'd254,  12'd0,  12'd42,  -12'd299,  
-12'd4,  -12'd140,  -12'd4,  -12'd32,  -12'd89,  12'd119,  -12'd98,  -12'd246,  12'd284,  12'd338,  -12'd337,  -12'd209,  -12'd199,  12'd381,  -12'd158,  -12'd596,  
-12'd73,  -12'd50,  -12'd327,  12'd60,  -12'd25,  -12'd158,  -12'd137,  -12'd24,  12'd247,  12'd154,  -12'd425,  12'd65,  -12'd184,  -12'd4,  -12'd207,  -12'd90,  
12'd114,  -12'd4,  -12'd119,  12'd120,  -12'd27,  12'd296,  -12'd426,  -12'd26,  12'd171,  -12'd53,  -12'd116,  -12'd321,  -12'd171,  -12'd156,  -12'd79,  -12'd313,  
12'd494,  -12'd140,  12'd180,  -12'd27,  -12'd931,  12'd352,  -12'd240,  -12'd42,  12'd81,  -12'd178,  -12'd196,  12'd607,  -12'd41,  12'd450,  12'd282,  -12'd177,  
12'd154,  -12'd96,  12'd262,  -12'd38,  -12'd33,  12'd224,  12'd586,  12'd219,  -12'd24,  12'd215,  12'd86,  12'd95,  12'd72,  12'd310,  12'd290,  -12'd105,  
12'd7,  -12'd248,  -12'd131,  -12'd120,  12'd152,  -12'd168,  12'd88,  12'd205,  12'd207,  -12'd368,  12'd114,  -12'd349,  -12'd134,  12'd22,  -12'd61,  12'd41,  
-12'd10,  -12'd136,  12'd191,  12'd263,  -12'd153,  -12'd221,  12'd73,  12'd31,  -12'd98,  -12'd139,  12'd33,  -12'd366,  12'd163,  -12'd38,  -12'd287,  -12'd105,  
-12'd370,  -12'd350,  -12'd240,  -12'd29,  12'd112,  -12'd222,  12'd40,  -12'd76,  12'd99,  12'd424,  -12'd248,  -12'd56,  12'd319,  -12'd199,  -12'd271,  12'd214,  

12'd201,  12'd272,  -12'd294,  -12'd246,  12'd318,  -12'd258,  -12'd312,  12'd445,  -12'd164,  12'd148,  12'd5,  12'd43,  12'd309,  12'd33,  -12'd326,  12'd301,  
-12'd157,  -12'd181,  -12'd238,  12'd163,  12'd303,  -12'd180,  -12'd512,  12'd333,  12'd57,  12'd36,  -12'd33,  12'd155,  12'd86,  12'd178,  12'd268,  12'd53,  
12'd294,  -12'd157,  -12'd76,  -12'd52,  -12'd310,  12'd282,  12'd160,  -12'd344,  12'd56,  -12'd317,  12'd578,  12'd32,  12'd163,  12'd179,  -12'd36,  12'd283,  
-12'd217,  -12'd183,  -12'd162,  12'd84,  -12'd53,  12'd6,  12'd511,  -12'd215,  -12'd215,  12'd59,  12'd101,  12'd91,  12'd252,  -12'd214,  12'd174,  -12'd118,  
-12'd89,  12'd39,  12'd16,  -12'd247,  -12'd283,  -12'd154,  12'd259,  12'd66,  -12'd170,  -12'd410,  12'd55,  -12'd228,  -12'd283,  12'd431,  12'd178,  12'd3,  
12'd7,  12'd39,  -12'd383,  -12'd29,  12'd58,  -12'd389,  -12'd438,  -12'd61,  -12'd155,  12'd132,  12'd416,  -12'd59,  -12'd73,  12'd43,  12'd37,  -12'd136,  
12'd315,  -12'd60,  12'd292,  12'd48,  12'd57,  -12'd221,  -12'd20,  -12'd355,  -12'd365,  12'd222,  12'd261,  12'd426,  12'd107,  -12'd110,  12'd154,  12'd172,  
-12'd136,  -12'd169,  12'd98,  12'd54,  12'd256,  -12'd479,  -12'd220,  12'd66,  -12'd249,  12'd483,  12'd475,  12'd272,  -12'd40,  -12'd1,  12'd219,  -12'd51,  
-12'd101,  -12'd19,  -12'd167,  -12'd292,  -12'd204,  -12'd542,  12'd129,  -12'd122,  -12'd231,  12'd373,  12'd8,  -12'd132,  12'd360,  -12'd9,  -12'd177,  12'd98,  
-12'd229,  12'd326,  12'd298,  -12'd365,  12'd72,  -12'd27,  -12'd53,  12'd402,  -12'd430,  12'd528,  -12'd161,  12'd263,  -12'd343,  12'd83,  -12'd434,  -12'd188,  
-12'd364,  -12'd338,  -12'd177,  -12'd322,  -12'd110,  12'd52,  -12'd253,  -12'd330,  12'd246,  12'd294,  12'd151,  -12'd42,  12'd74,  12'd144,  -12'd102,  12'd182,  
12'd49,  -12'd352,  -12'd94,  12'd265,  12'd62,  -12'd161,  -12'd515,  -12'd68,  12'd118,  12'd165,  -12'd111,  12'd26,  -12'd186,  12'd81,  -12'd356,  12'd301,  
12'd172,  -12'd401,  12'd48,  12'd258,  12'd111,  -12'd14,  12'd21,  12'd56,  12'd363,  12'd463,  -12'd257,  12'd128,  -12'd202,  -12'd308,  -12'd249,  12'd158,  
-12'd530,  12'd73,  -12'd98,  -12'd8,  12'd347,  -12'd79,  -12'd393,  12'd126,  12'd56,  12'd291,  -12'd237,  -12'd304,  12'd274,  -12'd101,  12'd306,  12'd312,  
-12'd165,  -12'd179,  -12'd372,  -12'd15,  12'd184,  12'd82,  -12'd51,  -12'd241,  12'd129,  12'd461,  -12'd36,  12'd324,  -12'd259,  12'd395,  12'd34,  -12'd319,  
-12'd197,  -12'd428,  12'd117,  -12'd101,  12'd172,  12'd19,  -12'd256,  -12'd211,  12'd452,  -12'd277,  12'd80,  -12'd278,  12'd234,  -12'd385,  12'd210,  12'd167,  
-12'd240,  -12'd288,  -12'd309,  -12'd74,  -12'd208,  12'd393,  -12'd389,  12'd205,  -12'd60,  12'd227,  12'd59,  12'd402,  12'd82,  -12'd255,  12'd86,  12'd53,  
12'd236,  -12'd157,  -12'd116,  12'd97,  -12'd199,  12'd350,  12'd112,  12'd318,  -12'd226,  -12'd263,  12'd333,  12'd248,  12'd5,  -12'd119,  -12'd6,  12'd17,  
-12'd3,  12'd400,  -12'd80,  12'd0,  12'd184,  -12'd15,  12'd57,  12'd325,  -12'd83,  12'd183,  -12'd58,  -12'd50,  -12'd100,  -12'd25,  -12'd44,  12'd56,  
-12'd20,  -12'd57,  12'd139,  -12'd13,  12'd412,  12'd53,  12'd51,  12'd437,  12'd290,  -12'd18,  12'd18,  -12'd375,  12'd77,  -12'd240,  12'd120,  12'd15,  
-12'd0,  -12'd142,  12'd200,  12'd276,  12'd90,  -12'd241,  12'd187,  -12'd93,  12'd155,  12'd97,  -12'd114,  12'd162,  12'd436,  12'd76,  12'd190,  12'd244,  
-12'd5,  -12'd102,  12'd12,  -12'd15,  -12'd327,  -12'd150,  12'd313,  12'd91,  12'd211,  -12'd463,  12'd144,  12'd108,  12'd265,  -12'd341,  12'd345,  12'd219,  
12'd364,  -12'd57,  -12'd293,  12'd135,  12'd153,  12'd95,  -12'd369,  -12'd21,  -12'd280,  12'd212,  12'd337,  12'd64,  12'd357,  -12'd230,  -12'd122,  -12'd215,  
12'd126,  12'd543,  -12'd124,  12'd290,  -12'd12,  -12'd121,  -12'd143,  12'd104,  12'd36,  -12'd24,  -12'd47,  12'd350,  12'd122,  -12'd253,  12'd1,  -12'd150,  
12'd506,  12'd363,  12'd199,  -12'd110,  -12'd32,  12'd143,  12'd89,  12'd46,  12'd498,  12'd796,  -12'd280,  12'd510,  12'd288,  12'd353,  12'd257,  12'd207,  

12'd334,  -12'd96,  -12'd428,  -12'd257,  12'd174,  -12'd31,  12'd178,  12'd136,  -12'd126,  12'd123,  12'd71,  -12'd157,  -12'd546,  12'd132,  12'd232,  -12'd114,  
-12'd292,  12'd10,  -12'd716,  12'd82,  12'd109,  12'd202,  12'd32,  -12'd38,  12'd223,  12'd53,  -12'd136,  12'd6,  -12'd374,  -12'd285,  -12'd176,  12'd111,  
-12'd29,  12'd77,  -12'd298,  12'd397,  -12'd144,  12'd410,  -12'd69,  -12'd40,  -12'd152,  12'd425,  12'd17,  12'd5,  12'd49,  -12'd478,  12'd246,  12'd44,  
-12'd232,  -12'd177,  -12'd162,  12'd209,  12'd53,  12'd31,  12'd24,  -12'd108,  12'd259,  12'd285,  -12'd113,  -12'd110,  12'd207,  -12'd254,  12'd53,  12'd303,  
-12'd173,  -12'd542,  -12'd136,  12'd213,  12'd194,  12'd64,  -12'd46,  12'd77,  -12'd40,  12'd256,  12'd65,  -12'd121,  -12'd436,  12'd182,  -12'd5,  12'd130,  
12'd218,  12'd153,  -12'd151,  -12'd141,  12'd18,  12'd66,  -12'd108,  12'd219,  12'd223,  12'd3,  12'd14,  12'd44,  12'd37,  12'd18,  12'd55,  12'd242,  
12'd329,  12'd311,  -12'd26,  -12'd312,  -12'd169,  -12'd3,  -12'd340,  -12'd18,  12'd245,  12'd146,  -12'd603,  -12'd168,  12'd78,  -12'd62,  12'd40,  12'd384,  
-12'd20,  -12'd86,  -12'd124,  -12'd146,  12'd149,  -12'd0,  12'd158,  -12'd117,  -12'd40,  12'd237,  12'd111,  12'd477,  -12'd69,  -12'd47,  12'd291,  12'd249,  
12'd131,  -12'd56,  -12'd697,  12'd312,  -12'd24,  12'd235,  -12'd109,  -12'd213,  12'd194,  12'd30,  -12'd219,  -12'd110,  -12'd58,  -12'd138,  12'd230,  12'd294,  
-12'd436,  -12'd373,  -12'd306,  12'd395,  -12'd404,  12'd15,  -12'd67,  12'd53,  12'd43,  -12'd589,  12'd141,  -12'd136,  12'd368,  12'd198,  -12'd97,  -12'd202,  
12'd43,  -12'd252,  12'd142,  12'd114,  12'd9,  -12'd211,  -12'd255,  12'd197,  12'd303,  12'd99,  -12'd504,  12'd172,  12'd459,  -12'd76,  12'd282,  12'd167,  
-12'd37,  -12'd140,  12'd199,  -12'd163,  -12'd251,  -12'd102,  12'd6,  12'd102,  -12'd8,  -12'd50,  -12'd290,  12'd42,  12'd193,  12'd381,  12'd49,  -12'd216,  
12'd322,  12'd69,  -12'd313,  12'd382,  12'd48,  -12'd56,  -12'd176,  12'd75,  -12'd138,  -12'd153,  12'd393,  -12'd6,  -12'd107,  -12'd171,  12'd139,  12'd111,  
12'd166,  12'd47,  12'd139,  12'd101,  -12'd379,  12'd265,  -12'd47,  12'd215,  -12'd123,  -12'd421,  12'd314,  12'd125,  12'd354,  12'd41,  -12'd241,  12'd285,  
-12'd93,  12'd293,  -12'd71,  12'd31,  12'd1,  12'd437,  12'd366,  12'd0,  12'd250,  12'd236,  12'd219,  -12'd231,  12'd78,  12'd275,  -12'd353,  12'd162,  
-12'd18,  -12'd143,  -12'd237,  -12'd80,  12'd503,  -12'd230,  -12'd350,  -12'd112,  -12'd117,  12'd259,  12'd331,  -12'd418,  -12'd15,  -12'd262,  12'd138,  -12'd182,  
-12'd257,  12'd283,  -12'd35,  -12'd52,  12'd105,  -12'd45,  -12'd444,  -12'd29,  -12'd69,  -12'd56,  -12'd264,  -12'd159,  -12'd37,  -12'd314,  -12'd252,  12'd251,  
12'd184,  -12'd189,  -12'd44,  -12'd88,  12'd60,  -12'd206,  12'd59,  -12'd1,  12'd217,  -12'd154,  12'd60,  12'd193,  -12'd458,  -12'd32,  -12'd16,  12'd224,  
12'd279,  12'd145,  -12'd181,  -12'd443,  -12'd177,  12'd53,  12'd166,  -12'd172,  -12'd102,  -12'd236,  12'd32,  12'd217,  -12'd227,  12'd133,  12'd52,  -12'd200,  
-12'd332,  12'd70,  -12'd256,  12'd218,  -12'd113,  -12'd221,  -12'd55,  12'd41,  -12'd203,  -12'd260,  12'd135,  -12'd170,  -12'd117,  12'd189,  12'd67,  -12'd271,  
-12'd79,  12'd132,  -12'd160,  -12'd130,  12'd384,  12'd364,  -12'd22,  -12'd120,  12'd448,  -12'd237,  12'd487,  12'd187,  12'd159,  -12'd323,  12'd328,  12'd240,  
-12'd123,  -12'd254,  -12'd240,  -12'd324,  12'd405,  -12'd328,  12'd57,  -12'd272,  -12'd53,  12'd142,  12'd52,  -12'd200,  -12'd113,  -12'd160,  -12'd85,  -12'd204,  
12'd87,  12'd231,  -12'd63,  -12'd154,  -12'd24,  -12'd98,  -12'd223,  -12'd525,  12'd456,  12'd347,  -12'd57,  12'd281,  -12'd163,  12'd494,  12'd30,  -12'd105,  
-12'd66,  12'd105,  -12'd8,  -12'd93,  -12'd194,  -12'd142,  -12'd22,  -12'd281,  12'd44,  -12'd55,  -12'd16,  12'd44,  12'd30,  12'd477,  -12'd216,  12'd61,  
-12'd375,  -12'd55,  12'd340,  12'd190,  12'd4,  -12'd57,  12'd115,  12'd221,  12'd304,  -12'd209,  -12'd96,  -12'd377,  -12'd346,  -12'd36,  -12'd34,  -12'd360,  

12'd205,  12'd195,  12'd325,  -12'd331,  -12'd85,  12'd176,  12'd204,  12'd50,  12'd329,  12'd18,  -12'd344,  -12'd143,  12'd75,  -12'd41,  -12'd112,  12'd142,  
-12'd275,  12'd472,  12'd292,  12'd138,  12'd379,  12'd33,  -12'd158,  -12'd122,  -12'd383,  -12'd76,  -12'd549,  12'd164,  12'd205,  -12'd142,  12'd183,  12'd173,  
12'd203,  -12'd159,  -12'd145,  12'd8,  -12'd194,  -12'd479,  12'd149,  -12'd125,  12'd114,  12'd53,  12'd6,  12'd157,  -12'd387,  12'd98,  12'd44,  12'd41,  
-12'd254,  -12'd327,  12'd390,  -12'd98,  -12'd114,  -12'd330,  -12'd76,  12'd82,  -12'd74,  -12'd288,  -12'd81,  -12'd230,  -12'd332,  12'd444,  12'd126,  12'd244,  
-12'd249,  12'd381,  12'd149,  12'd12,  -12'd189,  12'd99,  12'd96,  12'd27,  12'd373,  -12'd84,  -12'd49,  -12'd357,  -12'd268,  12'd411,  -12'd135,  12'd277,  
12'd63,  12'd193,  -12'd163,  -12'd193,  12'd180,  -12'd90,  12'd44,  12'd409,  -12'd181,  -12'd114,  -12'd323,  -12'd7,  -12'd419,  12'd85,  -12'd250,  12'd0,  
-12'd219,  -12'd150,  12'd49,  12'd51,  12'd343,  12'd117,  -12'd280,  12'd134,  -12'd86,  12'd212,  -12'd565,  12'd149,  -12'd178,  -12'd474,  12'd135,  -12'd218,  
-12'd123,  -12'd197,  12'd44,  -12'd115,  12'd10,  12'd179,  -12'd82,  -12'd273,  12'd88,  12'd258,  12'd11,  -12'd79,  -12'd185,  -12'd185,  -12'd139,  -12'd244,  
-12'd244,  -12'd436,  12'd355,  -12'd40,  -12'd137,  -12'd278,  -12'd6,  12'd61,  -12'd197,  -12'd94,  12'd168,  12'd45,  -12'd270,  12'd281,  12'd247,  -12'd229,  
-12'd258,  12'd54,  -12'd126,  -12'd107,  -12'd27,  12'd129,  -12'd31,  12'd499,  -12'd16,  12'd112,  -12'd107,  12'd80,  12'd158,  12'd219,  -12'd308,  -12'd537,  
12'd10,  -12'd70,  12'd80,  -12'd160,  12'd397,  -12'd0,  -12'd280,  12'd1,  12'd242,  12'd9,  -12'd360,  12'd95,  12'd268,  -12'd296,  -12'd239,  12'd10,  
12'd111,  12'd363,  12'd249,  12'd190,  -12'd250,  12'd217,  -12'd209,  12'd131,  -12'd203,  12'd333,  12'd378,  12'd178,  12'd240,  -12'd341,  12'd69,  12'd387,  
-12'd23,  -12'd265,  -12'd4,  12'd331,  12'd113,  12'd379,  -12'd169,  12'd481,  -12'd234,  -12'd188,  12'd462,  12'd224,  12'd306,  -12'd171,  -12'd150,  -12'd29,  
12'd31,  -12'd136,  -12'd111,  -12'd193,  -12'd226,  -12'd276,  12'd270,  -12'd352,  12'd353,  -12'd75,  12'd402,  -12'd18,  12'd110,  -12'd4,  -12'd193,  -12'd145,  
12'd166,  -12'd157,  -12'd540,  12'd272,  -12'd100,  12'd222,  12'd12,  12'd207,  12'd116,  -12'd179,  -12'd56,  12'd65,  12'd296,  -12'd253,  12'd191,  12'd265,  
12'd49,  -12'd357,  -12'd317,  12'd93,  12'd101,  12'd41,  12'd286,  12'd180,  12'd4,  12'd55,  12'd636,  12'd51,  12'd392,  12'd383,  12'd301,  12'd130,  
12'd254,  -12'd376,  12'd332,  12'd118,  12'd85,  12'd278,  12'd137,  -12'd63,  -12'd240,  12'd115,  -12'd40,  -12'd42,  12'd339,  12'd56,  12'd162,  12'd192,  
12'd7,  12'd365,  12'd365,  12'd272,  12'd75,  12'd127,  -12'd11,  -12'd209,  -12'd103,  -12'd73,  12'd345,  12'd15,  -12'd245,  -12'd211,  -12'd184,  12'd247,  
12'd31,  12'd183,  12'd72,  12'd60,  12'd468,  12'd50,  -12'd82,  -12'd15,  -12'd119,  -12'd116,  12'd145,  12'd30,  12'd72,  12'd46,  -12'd186,  -12'd223,  
12'd346,  -12'd73,  -12'd98,  12'd381,  -12'd353,  12'd211,  12'd40,  -12'd38,  12'd125,  12'd240,  -12'd21,  12'd82,  -12'd59,  12'd122,  -12'd33,  -12'd254,  
12'd219,  12'd252,  12'd276,  12'd76,  -12'd326,  -12'd33,  -12'd13,  -12'd6,  -12'd220,  12'd174,  12'd330,  -12'd280,  12'd348,  12'd237,  12'd108,  -12'd36,  
-12'd86,  12'd101,  -12'd217,  -12'd76,  -12'd41,  -12'd110,  12'd259,  -12'd73,  -12'd160,  -12'd47,  -12'd150,  -12'd27,  12'd377,  12'd142,  -12'd23,  -12'd90,  
12'd245,  12'd184,  12'd164,  12'd225,  -12'd1,  12'd182,  -12'd160,  -12'd195,  12'd258,  -12'd173,  12'd148,  -12'd135,  -12'd85,  -12'd94,  -12'd129,  -12'd37,  
-12'd348,  12'd398,  12'd228,  -12'd44,  -12'd215,  -12'd98,  -12'd173,  12'd236,  12'd225,  -12'd15,  -12'd179,  -12'd5,  -12'd73,  12'd240,  12'd237,  12'd423,  
12'd445,  12'd50,  12'd423,  12'd184,  12'd101,  -12'd62,  12'd209,  12'd265,  12'd317,  12'd66,  12'd134,  12'd386,  -12'd162,  12'd46,  12'd423,  12'd202,  

12'd19,  12'd103,  12'd475,  -12'd136,  -12'd465,  -12'd86,  12'd427,  -12'd213,  -12'd132,  -12'd403,  12'd115,  -12'd126,  -12'd286,  12'd447,  12'd207,  12'd28,  
-12'd179,  -12'd111,  12'd162,  -12'd2,  12'd257,  -12'd118,  12'd532,  -12'd508,  12'd189,  -12'd183,  12'd724,  -12'd145,  -12'd200,  12'd101,  -12'd263,  -12'd242,  
12'd90,  12'd39,  12'd27,  -12'd421,  -12'd10,  -12'd390,  -12'd32,  -12'd434,  12'd245,  12'd176,  12'd218,  12'd119,  12'd176,  12'd607,  -12'd175,  -12'd284,  
12'd240,  12'd225,  -12'd343,  -12'd72,  -12'd299,  -12'd137,  12'd185,  12'd159,  12'd305,  -12'd141,  12'd109,  -12'd326,  -12'd77,  -12'd337,  -12'd42,  -12'd163,  
12'd485,  12'd204,  -12'd194,  12'd459,  -12'd110,  12'd60,  -12'd240,  12'd174,  -12'd40,  -12'd77,  -12'd43,  12'd322,  12'd439,  12'd499,  12'd126,  12'd443,  
-12'd11,  12'd175,  12'd115,  -12'd226,  12'd5,  12'd110,  12'd407,  -12'd11,  -12'd370,  -12'd193,  -12'd191,  12'd304,  -12'd229,  12'd234,  -12'd96,  -12'd248,  
12'd196,  -12'd366,  -12'd89,  -12'd60,  -12'd42,  -12'd163,  12'd306,  12'd144,  12'd225,  -12'd326,  -12'd93,  12'd294,  12'd28,  12'd54,  12'd18,  -12'd129,  
-12'd32,  -12'd138,  12'd46,  12'd280,  12'd128,  -12'd37,  -12'd276,  -12'd451,  12'd311,  12'd595,  12'd328,  -12'd14,  -12'd233,  12'd144,  -12'd135,  -12'd203,  
-12'd42,  -12'd196,  -12'd769,  -12'd338,  -12'd24,  -12'd144,  -12'd412,  12'd180,  -12'd27,  12'd244,  12'd79,  -12'd469,  12'd323,  -12'd368,  -12'd233,  12'd128,  
-12'd388,  -12'd19,  -12'd201,  12'd97,  12'd271,  12'd312,  -12'd330,  -12'd77,  -12'd302,  12'd498,  12'd199,  12'd54,  12'd301,  -12'd253,  -12'd75,  12'd143,  
12'd37,  -12'd57,  12'd230,  12'd253,  -12'd156,  -12'd51,  12'd135,  -12'd125,  12'd244,  12'd92,  -12'd90,  12'd62,  12'd197,  12'd256,  12'd419,  12'd232,  
12'd104,  -12'd213,  12'd351,  12'd456,  -12'd136,  12'd111,  -12'd215,  12'd488,  -12'd51,  12'd88,  12'd23,  -12'd212,  12'd440,  12'd393,  12'd286,  -12'd275,  
-12'd103,  -12'd306,  -12'd114,  12'd176,  12'd405,  12'd37,  12'd125,  -12'd352,  -12'd17,  12'd45,  12'd270,  12'd127,  12'd88,  -12'd359,  12'd13,  -12'd241,  
-12'd166,  -12'd146,  -12'd649,  -12'd90,  -12'd17,  12'd143,  -12'd188,  -12'd99,  12'd259,  -12'd315,  12'd191,  12'd21,  12'd87,  -12'd349,  -12'd238,  -12'd125,  
-12'd432,  12'd3,  -12'd141,  12'd523,  -12'd48,  12'd123,  -12'd465,  12'd196,  12'd57,  12'd265,  12'd444,  -12'd172,  12'd143,  -12'd41,  12'd108,  -12'd142,  
12'd55,  12'd35,  12'd178,  12'd2,  -12'd9,  12'd222,  12'd88,  -12'd159,  -12'd244,  -12'd10,  -12'd33,  12'd67,  12'd192,  12'd78,  -12'd88,  -12'd61,  
12'd8,  -12'd169,  12'd39,  12'd258,  12'd255,  -12'd323,  -12'd600,  -12'd94,  -12'd320,  -12'd50,  -12'd144,  12'd95,  12'd83,  12'd86,  12'd98,  12'd150,  
12'd328,  12'd61,  12'd466,  -12'd40,  12'd177,  12'd10,  12'd316,  -12'd139,  -12'd198,  12'd47,  -12'd54,  12'd418,  12'd314,  12'd238,  12'd1,  12'd72,  
12'd64,  -12'd19,  12'd18,  -12'd110,  12'd560,  12'd24,  12'd50,  -12'd86,  12'd166,  -12'd241,  12'd410,  12'd261,  -12'd113,  12'd126,  -12'd28,  -12'd110,  
-12'd1,  12'd189,  12'd99,  -12'd46,  12'd176,  12'd48,  12'd11,  12'd242,  12'd69,  -12'd102,  -12'd187,  -12'd230,  -12'd428,  12'd207,  -12'd31,  -12'd278,  
12'd292,  12'd49,  -12'd120,  -12'd150,  -12'd62,  12'd32,  12'd332,  12'd31,  12'd276,  12'd72,  -12'd45,  12'd25,  12'd120,  -12'd69,  -12'd200,  12'd138,  
-12'd183,  -12'd156,  12'd19,  -12'd50,  -12'd178,  -12'd105,  -12'd191,  -12'd229,  12'd239,  12'd125,  12'd355,  -12'd43,  12'd198,  -12'd586,  12'd197,  12'd179,  
-12'd192,  12'd90,  12'd261,  12'd48,  -12'd200,  -12'd402,  12'd135,  -12'd64,  12'd220,  12'd232,  12'd95,  12'd63,  -12'd87,  12'd338,  12'd12,  12'd85,  
-12'd264,  12'd58,  12'd309,  -12'd169,  -12'd250,  -12'd100,  -12'd67,  12'd235,  12'd139,  -12'd179,  -12'd352,  -12'd43,  12'd214,  12'd61,  12'd124,  -12'd113,  
-12'd182,  12'd93,  12'd3,  -12'd29,  -12'd338,  12'd99,  -12'd165,  12'd235,  -12'd162,  -12'd377,  -12'd184,  -12'd312,  -12'd12,  12'd370,  12'd193,  -12'd331,  

-12'd0,  12'd169,  -12'd120,  12'd62,  -12'd380,  -12'd137,  12'd256,  12'd157,  12'd195,  12'd8,  -12'd132,  -12'd25,  -12'd127,  -12'd166,  12'd431,  12'd73,  
-12'd40,  12'd157,  -12'd23,  12'd153,  -12'd19,  12'd220,  -12'd174,  12'd245,  12'd204,  12'd204,  12'd446,  -12'd226,  -12'd340,  -12'd474,  12'd115,  12'd96,  
12'd175,  12'd152,  -12'd179,  12'd129,  12'd87,  12'd131,  -12'd546,  -12'd0,  12'd57,  12'd12,  12'd343,  -12'd32,  12'd258,  -12'd659,  12'd80,  -12'd85,  
12'd16,  -12'd141,  12'd178,  -12'd15,  -12'd210,  12'd182,  -12'd431,  12'd172,  -12'd43,  12'd72,  -12'd162,  -12'd27,  12'd43,  -12'd947,  -12'd34,  12'd143,  
-12'd344,  -12'd394,  12'd79,  -12'd214,  -12'd100,  -12'd211,  -12'd245,  -12'd25,  12'd138,  12'd133,  -12'd81,  12'd186,  -12'd163,  12'd75,  -12'd163,  12'd7,  
-12'd17,  -12'd243,  12'd524,  12'd426,  -12'd92,  12'd125,  -12'd194,  12'd175,  -12'd52,  -12'd16,  12'd65,  12'd170,  12'd201,  -12'd175,  12'd9,  12'd110,  
-12'd384,  -12'd179,  -12'd74,  -12'd33,  12'd150,  12'd278,  12'd287,  12'd120,  12'd114,  -12'd48,  -12'd72,  12'd52,  -12'd200,  -12'd211,  -12'd29,  12'd84,  
-12'd542,  -12'd64,  -12'd379,  12'd359,  12'd175,  12'd252,  -12'd427,  -12'd120,  -12'd186,  -12'd53,  -12'd123,  -12'd225,  -12'd235,  -12'd368,  -12'd80,  -12'd231,  
-12'd290,  12'd234,  12'd0,  -12'd302,  12'd254,  12'd21,  -12'd217,  -12'd302,  -12'd361,  12'd380,  -12'd215,  -12'd332,  -12'd111,  -12'd160,  12'd49,  12'd154,  
-12'd637,  -12'd54,  12'd68,  -12'd44,  -12'd177,  -12'd178,  12'd134,  12'd33,  12'd102,  12'd190,  12'd84,  -12'd454,  -12'd135,  12'd39,  -12'd69,  -12'd306,  
12'd46,  12'd83,  12'd176,  12'd258,  12'd210,  12'd107,  -12'd34,  12'd232,  -12'd468,  12'd2,  12'd162,  12'd241,  12'd264,  12'd225,  12'd105,  12'd88,  
-12'd368,  12'd163,  -12'd199,  12'd57,  12'd435,  -12'd52,  -12'd123,  12'd42,  12'd473,  12'd79,  12'd246,  12'd223,  12'd49,  -12'd493,  -12'd58,  -12'd98,  
12'd71,  12'd150,  12'd28,  -12'd109,  12'd427,  12'd29,  12'd9,  12'd91,  12'd5,  12'd119,  12'd94,  12'd208,  -12'd306,  12'd193,  -12'd176,  12'd308,  
12'd186,  -12'd350,  12'd349,  -12'd58,  -12'd295,  -12'd66,  -12'd76,  -12'd21,  -12'd217,  -12'd462,  12'd185,  -12'd24,  12'd60,  12'd212,  12'd250,  -12'd81,  
12'd281,  -12'd297,  12'd352,  -12'd261,  -12'd67,  12'd413,  -12'd77,  12'd77,  12'd265,  12'd80,  -12'd41,  -12'd60,  12'd31,  12'd229,  -12'd6,  12'd164,  
12'd511,  12'd12,  12'd51,  -12'd290,  -12'd263,  -12'd141,  12'd217,  -12'd218,  12'd300,  -12'd23,  12'd249,  12'd378,  -12'd286,  -12'd307,  12'd7,  -12'd229,  
-12'd19,  -12'd82,  -12'd385,  12'd104,  -12'd49,  -12'd92,  -12'd40,  -12'd270,  12'd452,  -12'd135,  12'd22,  12'd373,  12'd223,  12'd165,  -12'd307,  12'd299,  
12'd186,  -12'd168,  -12'd86,  12'd7,  -12'd220,  12'd276,  12'd271,  -12'd146,  12'd150,  -12'd97,  -12'd266,  12'd83,  12'd215,  -12'd137,  -12'd189,  12'd122,  
12'd291,  12'd172,  12'd383,  12'd196,  12'd267,  -12'd179,  12'd37,  12'd116,  -12'd22,  -12'd107,  12'd125,  -12'd393,  12'd198,  12'd0,  12'd199,  12'd13,  
-12'd291,  12'd328,  -12'd237,  -12'd71,  -12'd60,  -12'd316,  -12'd218,  -12'd66,  -12'd127,  12'd476,  12'd75,  12'd55,  12'd371,  -12'd41,  12'd113,  -12'd208,  
12'd359,  12'd304,  12'd85,  -12'd89,  12'd108,  -12'd11,  12'd638,  -12'd93,  -12'd118,  -12'd394,  12'd81,  12'd304,  -12'd251,  -12'd124,  -12'd354,  12'd150,  
12'd28,  12'd101,  -12'd351,  -12'd133,  -12'd122,  -12'd67,  12'd707,  -12'd142,  12'd386,  12'd145,  12'd150,  -12'd99,  -12'd151,  12'd283,  -12'd363,  -12'd312,  
12'd59,  -12'd136,  12'd226,  -12'd73,  12'd8,  -12'd162,  -12'd51,  -12'd81,  12'd140,  12'd27,  -12'd31,  -12'd360,  12'd228,  12'd340,  -12'd142,  -12'd280,  
-12'd30,  12'd376,  12'd45,  -12'd123,  -12'd97,  12'd455,  -12'd83,  12'd110,  -12'd30,  12'd203,  12'd79,  -12'd172,  12'd118,  -12'd199,  12'd18,  12'd96,  
-12'd546,  -12'd465,  -12'd438,  12'd321,  12'd61,  12'd282,  12'd134,  -12'd140,  -12'd202,  12'd340,  -12'd238,  -12'd383,  -12'd171,  -12'd387,  12'd272,  -12'd118,  

12'd293,  12'd93,  12'd26,  12'd48,  -12'd156,  12'd93,  12'd440,  12'd107,  12'd109,  -12'd104,  12'd219,  12'd152,  12'd22,  12'd184,  -12'd30,  12'd119,  
12'd128,  12'd184,  12'd319,  12'd161,  12'd173,  12'd105,  12'd61,  -12'd16,  12'd231,  12'd212,  12'd514,  12'd63,  12'd72,  12'd269,  -12'd11,  -12'd184,  
-12'd179,  -12'd407,  12'd173,  -12'd49,  12'd49,  12'd234,  12'd351,  12'd372,  -12'd67,  12'd249,  12'd212,  12'd176,  12'd85,  -12'd165,  12'd216,  12'd160,  
-12'd54,  -12'd211,  12'd185,  12'd147,  -12'd281,  -12'd48,  -12'd56,  -12'd51,  -12'd124,  12'd305,  -12'd311,  -12'd18,  12'd275,  -12'd92,  -12'd185,  12'd2,  
-12'd154,  -12'd135,  -12'd321,  -12'd279,  -12'd12,  -12'd195,  -12'd39,  -12'd17,  -12'd158,  12'd41,  12'd8,  -12'd177,  12'd177,  12'd58,  -12'd119,  -12'd132,  
-12'd10,  12'd246,  -12'd105,  12'd186,  12'd110,  12'd289,  -12'd127,  -12'd32,  12'd135,  12'd220,  -12'd32,  -12'd189,  -12'd251,  12'd325,  12'd37,  -12'd277,  
-12'd94,  12'd22,  12'd281,  -12'd254,  -12'd162,  -12'd313,  -12'd22,  12'd45,  12'd112,  12'd39,  12'd257,  12'd28,  -12'd34,  12'd326,  12'd49,  12'd243,  
-12'd36,  -12'd349,  12'd14,  12'd138,  -12'd60,  12'd210,  -12'd27,  12'd111,  12'd4,  12'd94,  -12'd298,  -12'd132,  12'd267,  12'd210,  12'd83,  12'd108,  
-12'd121,  -12'd449,  12'd1,  12'd175,  12'd201,  12'd136,  -12'd48,  12'd120,  -12'd66,  -12'd184,  -12'd134,  -12'd298,  -12'd64,  12'd25,  -12'd52,  12'd11,  
-12'd808,  -12'd294,  -12'd404,  -12'd162,  -12'd274,  -12'd591,  -12'd29,  -12'd81,  -12'd497,  -12'd52,  -12'd26,  12'd144,  -12'd436,  12'd158,  -12'd234,  -12'd132,  
-12'd357,  -12'd392,  12'd371,  -12'd77,  12'd136,  12'd145,  -12'd190,  12'd293,  12'd171,  12'd344,  -12'd366,  -12'd66,  12'd24,  12'd572,  12'd255,  -12'd51,  
12'd15,  -12'd110,  12'd176,  12'd244,  -12'd51,  -12'd96,  -12'd336,  -12'd47,  -12'd353,  -12'd415,  -12'd34,  12'd4,  12'd114,  12'd15,  12'd393,  12'd95,  
12'd23,  -12'd98,  12'd241,  12'd201,  -12'd303,  12'd129,  -12'd488,  -12'd181,  12'd188,  12'd150,  -12'd111,  -12'd240,  12'd27,  -12'd238,  12'd51,  -12'd33,  
12'd96,  -12'd208,  -12'd83,  -12'd172,  -12'd58,  12'd166,  -12'd193,  -12'd225,  -12'd254,  -12'd154,  -12'd289,  -12'd135,  -12'd247,  12'd118,  12'd49,  -12'd370,  
-12'd3,  -12'd144,  12'd35,  12'd33,  -12'd317,  12'd75,  12'd65,  12'd74,  12'd75,  12'd304,  -12'd140,  12'd51,  -12'd410,  -12'd146,  -12'd316,  12'd98,  
-12'd408,  12'd115,  -12'd147,  -12'd54,  12'd352,  12'd115,  -12'd346,  12'd339,  12'd28,  12'd346,  -12'd370,  -12'd33,  12'd37,  12'd60,  -12'd298,  -12'd216,  
-12'd241,  12'd339,  12'd163,  -12'd67,  -12'd295,  12'd26,  -12'd534,  12'd14,  12'd132,  -12'd121,  12'd255,  12'd61,  -12'd275,  -12'd200,  -12'd75,  -12'd94,  
-12'd329,  -12'd84,  12'd37,  -12'd323,  12'd16,  -12'd423,  12'd209,  12'd108,  -12'd432,  -12'd79,  -12'd145,  12'd234,  12'd118,  12'd31,  -12'd90,  12'd346,  
12'd87,  12'd89,  12'd19,  12'd60,  -12'd295,  -12'd144,  12'd18,  12'd11,  12'd303,  12'd44,  -12'd112,  12'd412,  12'd28,  12'd254,  12'd383,  -12'd86,  
-12'd221,  12'd107,  12'd176,  -12'd392,  -12'd342,  12'd145,  12'd352,  12'd146,  -12'd280,  12'd323,  12'd3,  12'd7,  -12'd160,  -12'd180,  12'd216,  -12'd406,  
-12'd499,  12'd94,  -12'd413,  12'd126,  12'd422,  -12'd306,  12'd223,  -12'd145,  12'd535,  -12'd75,  -12'd8,  -12'd165,  -12'd163,  -12'd156,  -12'd91,  -12'd116,  
-12'd11,  -12'd112,  -12'd340,  -12'd77,  12'd448,  12'd219,  12'd86,  -12'd468,  12'd165,  12'd123,  12'd279,  12'd27,  -12'd156,  -12'd406,  -12'd9,  12'd270,  
12'd256,  12'd278,  -12'd82,  12'd0,  -12'd137,  -12'd172,  -12'd86,  -12'd158,  12'd250,  12'd80,  12'd124,  12'd218,  12'd105,  12'd166,  -12'd78,  -12'd237,  
12'd306,  12'd172,  12'd214,  12'd123,  12'd295,  12'd513,  12'd183,  12'd243,  -12'd114,  12'd86,  -12'd43,  12'd247,  12'd414,  -12'd3,  12'd5,  12'd193,  
12'd212,  -12'd144,  12'd378,  -12'd6,  12'd83,  12'd157,  12'd311,  12'd243,  12'd77,  -12'd299,  -12'd3,  12'd375,  12'd83,  12'd2,  12'd31,  -12'd86,  

12'd430,  12'd39,  12'd453,  12'd134,  12'd7,  12'd223,  12'd87,  -12'd421,  -12'd88,  12'd135,  12'd152,  12'd151,  -12'd71,  -12'd190,  12'd69,  -12'd37,  
-12'd22,  12'd204,  12'd389,  -12'd7,  -12'd6,  12'd182,  -12'd69,  -12'd114,  12'd20,  -12'd194,  -12'd195,  12'd98,  -12'd91,  -12'd66,  -12'd2,  12'd148,  
12'd50,  12'd43,  -12'd324,  12'd136,  12'd77,  12'd31,  12'd69,  12'd216,  12'd255,  -12'd113,  12'd68,  12'd19,  -12'd324,  12'd93,  -12'd178,  12'd148,  
12'd41,  -12'd155,  12'd147,  -12'd474,  12'd67,  -12'd41,  12'd92,  -12'd120,  12'd338,  12'd34,  12'd69,  12'd349,  -12'd327,  12'd755,  -12'd261,  -12'd263,  
-12'd103,  12'd80,  12'd274,  12'd173,  12'd8,  12'd71,  12'd76,  -12'd14,  12'd208,  -12'd31,  -12'd23,  -12'd69,  -12'd207,  12'd483,  -12'd236,  -12'd134,  
-12'd61,  12'd315,  -12'd183,  -12'd150,  -12'd130,  12'd332,  12'd154,  -12'd69,  -12'd54,  12'd7,  12'd39,  -12'd57,  -12'd154,  12'd64,  12'd80,  12'd27,  
-12'd11,  -12'd80,  12'd341,  -12'd315,  -12'd54,  12'd286,  12'd73,  12'd211,  -12'd145,  12'd10,  -12'd239,  -12'd12,  -12'd134,  12'd223,  12'd477,  -12'd133,  
12'd605,  -12'd292,  12'd415,  12'd190,  12'd189,  12'd9,  12'd366,  -12'd60,  -12'd50,  12'd35,  -12'd101,  12'd282,  -12'd110,  -12'd2,  12'd91,  -12'd411,  
-12'd39,  -12'd308,  -12'd34,  12'd237,  12'd153,  12'd18,  12'd138,  -12'd334,  12'd64,  -12'd104,  -12'd411,  12'd9,  12'd305,  12'd386,  -12'd197,  -12'd103,  
12'd91,  -12'd28,  -12'd180,  12'd177,  12'd456,  12'd314,  12'd269,  12'd87,  12'd190,  -12'd164,  -12'd219,  -12'd241,  12'd51,  12'd382,  -12'd509,  -12'd167,  
-12'd82,  12'd379,  12'd2,  12'd56,  12'd28,  -12'd94,  12'd343,  12'd82,  -12'd176,  -12'd133,  12'd16,  -12'd258,  12'd113,  -12'd87,  -12'd190,  12'd253,  
-12'd105,  -12'd180,  12'd163,  12'd239,  12'd384,  12'd367,  12'd278,  12'd178,  12'd120,  -12'd275,  -12'd335,  -12'd301,  12'd214,  12'd254,  -12'd233,  12'd12,  
12'd333,  12'd204,  -12'd108,  -12'd25,  -12'd17,  12'd423,  -12'd193,  12'd96,  12'd212,  -12'd333,  -12'd187,  12'd96,  12'd174,  -12'd402,  12'd418,  -12'd335,  
12'd32,  -12'd39,  12'd69,  -12'd122,  -12'd3,  12'd44,  12'd76,  -12'd229,  -12'd157,  12'd80,  -12'd74,  12'd33,  -12'd16,  12'd106,  12'd259,  12'd173,  
12'd160,  -12'd475,  -12'd177,  -12'd89,  12'd366,  12'd147,  12'd346,  12'd107,  -12'd152,  12'd147,  -12'd294,  -12'd254,  -12'd41,  12'd476,  12'd49,  12'd92,  
12'd287,  12'd187,  12'd170,  12'd201,  -12'd326,  -12'd111,  12'd208,  12'd145,  12'd66,  -12'd9,  -12'd14,  -12'd14,  -12'd44,  12'd198,  -12'd144,  12'd160,  
12'd292,  -12'd70,  12'd48,  12'd130,  12'd626,  -12'd88,  12'd179,  12'd132,  12'd314,  12'd11,  -12'd188,  -12'd155,  -12'd10,  12'd452,  -12'd95,  12'd56,  
12'd55,  12'd104,  -12'd51,  12'd16,  12'd175,  12'd16,  -12'd161,  -12'd229,  -12'd119,  -12'd216,  -12'd372,  12'd56,  -12'd330,  12'd341,  -12'd21,  12'd177,  
-12'd0,  -12'd399,  12'd205,  -12'd176,  -12'd136,  12'd57,  12'd10,  12'd67,  12'd265,  -12'd335,  -12'd229,  12'd157,  -12'd157,  -12'd61,  12'd150,  12'd96,  
-12'd326,  12'd26,  -12'd16,  12'd24,  -12'd220,  12'd4,  12'd466,  12'd5,  12'd306,  -12'd382,  -12'd39,  -12'd136,  -12'd30,  -12'd305,  -12'd2,  12'd87,  
12'd127,  12'd31,  -12'd68,  12'd175,  -12'd9,  -12'd344,  -12'd371,  -12'd60,  -12'd314,  12'd148,  -12'd509,  -12'd322,  12'd2,  12'd294,  -12'd30,  12'd91,  
-12'd134,  12'd385,  12'd65,  12'd140,  12'd181,  -12'd100,  -12'd213,  12'd55,  -12'd277,  12'd11,  -12'd389,  -12'd191,  -12'd64,  12'd335,  12'd299,  12'd56,  
12'd233,  12'd269,  12'd92,  -12'd288,  -12'd45,  12'd50,  12'd17,  12'd230,  -12'd6,  -12'd246,  -12'd261,  -12'd260,  -12'd231,  12'd437,  12'd597,  -12'd172,  
12'd132,  -12'd212,  12'd114,  12'd23,  12'd284,  -12'd188,  12'd298,  12'd302,  -12'd136,  -12'd467,  -12'd170,  -12'd248,  12'd147,  12'd554,  12'd190,  12'd351,  
12'd43,  12'd285,  -12'd30,  12'd206,  12'd529,  12'd364,  12'd135,  12'd168,  -12'd158,  -12'd456,  12'd47,  -12'd82,  -12'd189,  12'd256,  12'd28,  -12'd265,  

12'd242,  -12'd252,  -12'd433,  12'd14,  -12'd101,  12'd16,  -12'd290,  -12'd17,  -12'd21,  12'd241,  -12'd446,  -12'd14,  12'd326,  12'd58,  12'd420,  12'd139,  
-12'd43,  12'd116,  12'd171,  12'd109,  -12'd94,  12'd12,  -12'd509,  12'd519,  12'd222,  12'd350,  12'd52,  -12'd60,  -12'd84,  -12'd39,  12'd240,  12'd127,  
-12'd3,  -12'd353,  12'd251,  12'd77,  -12'd238,  12'd34,  -12'd46,  12'd264,  12'd109,  12'd29,  12'd0,  12'd272,  -12'd96,  -12'd120,  12'd276,  12'd59,  
12'd90,  12'd84,  12'd413,  12'd96,  -12'd403,  -12'd290,  -12'd441,  12'd18,  12'd37,  12'd219,  -12'd178,  12'd161,  12'd293,  -12'd419,  12'd235,  -12'd268,  
12'd180,  12'd296,  12'd60,  12'd256,  -12'd207,  -12'd96,  12'd55,  12'd300,  12'd48,  12'd197,  -12'd11,  12'd53,  12'd259,  -12'd317,  12'd82,  12'd287,  
12'd24,  12'd280,  -12'd58,  12'd403,  12'd54,  12'd243,  -12'd504,  -12'd268,  12'd285,  12'd420,  -12'd324,  12'd54,  12'd250,  -12'd178,  12'd172,  -12'd274,  
-12'd234,  12'd38,  12'd155,  12'd342,  -12'd143,  12'd28,  -12'd90,  12'd0,  12'd119,  12'd399,  -12'd192,  -12'd245,  12'd214,  12'd411,  12'd165,  12'd73,  
12'd8,  12'd245,  12'd446,  12'd181,  12'd85,  -12'd352,  12'd27,  -12'd192,  12'd150,  -12'd28,  12'd292,  -12'd58,  12'd233,  12'd481,  -12'd153,  12'd372,  
-12'd242,  12'd345,  12'd168,  -12'd109,  -12'd145,  12'd226,  -12'd59,  12'd131,  -12'd253,  -12'd108,  12'd206,  12'd169,  -12'd53,  12'd89,  12'd70,  -12'd194,  
12'd338,  -12'd180,  12'd145,  12'd59,  -12'd315,  12'd238,  12'd120,  12'd161,  -12'd101,  -12'd162,  12'd53,  12'd425,  12'd101,  -12'd320,  -12'd141,  -12'd282,  
-12'd232,  12'd255,  -12'd16,  12'd31,  12'd300,  -12'd50,  -12'd463,  12'd372,  -12'd384,  -12'd88,  -12'd97,  12'd57,  -12'd215,  12'd88,  12'd18,  -12'd6,  
12'd24,  12'd157,  12'd77,  -12'd101,  12'd373,  12'd16,  12'd358,  -12'd53,  12'd67,  12'd141,  12'd87,  12'd58,  12'd7,  -12'd279,  -12'd125,  12'd52,  
-12'd239,  -12'd363,  12'd333,  -12'd283,  12'd234,  12'd221,  12'd143,  12'd80,  12'd56,  12'd89,  12'd161,  12'd170,  -12'd420,  12'd499,  12'd18,  -12'd307,  
12'd112,  -12'd191,  -12'd152,  12'd362,  12'd169,  -12'd408,  -12'd48,  12'd334,  12'd88,  12'd20,  -12'd128,  -12'd168,  -12'd0,  -12'd72,  12'd112,  -12'd27,  
12'd467,  12'd386,  12'd5,  -12'd231,  12'd14,  -12'd289,  -12'd50,  12'd144,  -12'd46,  -12'd407,  -12'd252,  -12'd96,  -12'd45,  12'd42,  12'd363,  12'd210,  
12'd170,  -12'd177,  -12'd96,  -12'd143,  -12'd88,  -12'd477,  12'd151,  -12'd322,  12'd124,  -12'd112,  -12'd239,  12'd465,  12'd96,  -12'd207,  -12'd190,  -12'd19,  
12'd397,  12'd178,  12'd68,  -12'd17,  -12'd74,  12'd68,  12'd905,  -12'd150,  12'd620,  -12'd24,  12'd145,  12'd18,  12'd208,  12'd474,  -12'd31,  12'd135,  
-12'd214,  12'd90,  -12'd58,  12'd63,  12'd75,  12'd276,  -12'd44,  -12'd194,  12'd238,  -12'd262,  12'd125,  -12'd152,  -12'd10,  12'd33,  -12'd176,  12'd104,  
-12'd365,  -12'd45,  -12'd209,  12'd106,  -12'd55,  -12'd279,  12'd162,  -12'd462,  12'd80,  12'd397,  -12'd193,  -12'd453,  -12'd256,  -12'd236,  -12'd35,  -12'd335,  
-12'd197,  12'd12,  -12'd49,  -12'd45,  12'd75,  -12'd144,  12'd42,  -12'd59,  -12'd131,  12'd356,  -12'd34,  12'd48,  -12'd205,  -12'd365,  12'd37,  12'd306,  
12'd99,  -12'd86,  12'd453,  -12'd122,  -12'd154,  -12'd107,  12'd365,  12'd14,  12'd84,  12'd142,  -12'd3,  -12'd190,  12'd249,  12'd506,  -12'd183,  12'd140,  
-12'd43,  12'd51,  12'd169,  12'd159,  -12'd103,  12'd93,  -12'd214,  12'd212,  -12'd489,  -12'd186,  -12'd135,  -12'd35,  -12'd12,  12'd421,  -12'd26,  12'd50,  
12'd311,  -12'd299,  -12'd227,  -12'd299,  -12'd326,  -12'd280,  -12'd395,  12'd56,  -12'd452,  -12'd337,  12'd205,  -12'd89,  -12'd79,  -12'd12,  12'd86,  12'd335,  
12'd404,  12'd127,  -12'd252,  -12'd40,  -12'd406,  -12'd120,  -12'd227,  12'd174,  -12'd95,  -12'd117,  12'd37,  -12'd51,  12'd173,  12'd135,  12'd18,  12'd157,  
12'd5,  12'd264,  12'd517,  -12'd355,  12'd61,  -12'd79,  12'd124,  -12'd1,  -12'd74,  -12'd454,  -12'd82,  -12'd54,  -12'd67,  -12'd105,  -12'd160,  12'd110,  

-12'd121,  -12'd455,  -12'd118,  12'd219,  12'd424,  -12'd126,  -12'd467,  -12'd170,  12'd5,  12'd283,  -12'd372,  12'd229,  12'd120,  -12'd423,  12'd164,  -12'd272,  
12'd308,  -12'd362,  -12'd124,  -12'd84,  12'd396,  12'd12,  -12'd112,  12'd19,  -12'd192,  12'd37,  -12'd150,  -12'd36,  12'd131,  12'd153,  12'd164,  -12'd194,  
12'd195,  -12'd41,  12'd393,  12'd106,  -12'd205,  -12'd55,  -12'd47,  12'd3,  12'd82,  -12'd156,  -12'd219,  12'd422,  -12'd277,  12'd53,  12'd249,  -12'd176,  
12'd115,  12'd30,  12'd265,  12'd240,  -12'd86,  12'd71,  12'd114,  12'd291,  -12'd167,  -12'd220,  -12'd28,  12'd102,  -12'd97,  12'd0,  12'd214,  -12'd139,  
12'd334,  12'd52,  12'd141,  12'd546,  -12'd28,  12'd42,  -12'd25,  -12'd198,  12'd344,  -12'd68,  -12'd109,  12'd133,  -12'd20,  -12'd484,  12'd407,  -12'd224,  
-12'd33,  12'd38,  12'd167,  12'd460,  -12'd303,  12'd327,  12'd58,  -12'd132,  -12'd54,  12'd0,  -12'd229,  12'd320,  -12'd221,  12'd241,  12'd17,  -12'd40,  
12'd223,  -12'd463,  -12'd341,  12'd52,  -12'd217,  12'd233,  12'd35,  12'd210,  12'd192,  12'd169,  12'd32,  12'd14,  -12'd80,  -12'd138,  12'd172,  12'd261,  
-12'd137,  -12'd167,  -12'd73,  12'd265,  -12'd45,  -12'd164,  12'd13,  12'd29,  -12'd205,  12'd14,  -12'd285,  -12'd25,  -12'd194,  12'd551,  12'd43,  -12'd75,  
12'd62,  12'd44,  -12'd48,  -12'd144,  -12'd41,  -12'd53,  -12'd187,  12'd482,  -12'd501,  -12'd333,  -12'd251,  12'd104,  12'd19,  12'd90,  12'd482,  -12'd86,  
12'd452,  12'd591,  12'd451,  -12'd176,  -12'd313,  -12'd24,  12'd69,  -12'd202,  12'd63,  -12'd498,  -12'd174,  12'd45,  -12'd448,  -12'd3,  12'd465,  12'd106,  
-12'd173,  12'd288,  12'd292,  12'd68,  12'd73,  -12'd15,  12'd504,  -12'd62,  12'd336,  12'd134,  -12'd158,  -12'd233,  -12'd74,  -12'd78,  12'd179,  12'd121,  
12'd27,  -12'd437,  -12'd156,  -12'd241,  12'd324,  -12'd186,  12'd490,  -12'd131,  -12'd10,  -12'd241,  -12'd78,  12'd239,  12'd297,  12'd384,  12'd41,  12'd34,  
-12'd369,  12'd256,  12'd104,  -12'd160,  -12'd162,  -12'd336,  -12'd182,  12'd464,  -12'd540,  12'd170,  -12'd26,  -12'd166,  -12'd212,  12'd126,  12'd136,  -12'd15,  
-12'd118,  -12'd17,  12'd426,  -12'd216,  -12'd320,  12'd21,  -12'd182,  12'd421,  12'd59,  -12'd435,  -12'd22,  12'd126,  -12'd494,  12'd45,  12'd404,  -12'd52,  
12'd54,  -12'd4,  12'd455,  12'd60,  -12'd270,  -12'd220,  -12'd191,  12'd261,  12'd44,  -12'd303,  -12'd351,  12'd159,  -12'd285,  -12'd153,  12'd94,  -12'd111,  
12'd3,  12'd48,  -12'd163,  -12'd25,  -12'd56,  12'd282,  12'd471,  12'd134,  -12'd313,  -12'd60,  -12'd50,  -12'd207,  12'd54,  -12'd89,  12'd169,  12'd301,  
12'd141,  -12'd19,  12'd39,  12'd374,  12'd295,  -12'd66,  -12'd84,  12'd237,  -12'd164,  -12'd260,  -12'd211,  -12'd205,  12'd92,  -12'd350,  12'd88,  -12'd279,  
-12'd279,  12'd37,  -12'd57,  -12'd212,  -12'd80,  -12'd438,  -12'd209,  12'd222,  -12'd351,  12'd249,  -12'd9,  -12'd436,  12'd57,  12'd284,  12'd4,  -12'd382,  
12'd18,  12'd12,  12'd383,  12'd41,  12'd186,  12'd233,  12'd283,  -12'd163,  12'd116,  -12'd287,  12'd91,  12'd341,  12'd64,  -12'd171,  -12'd207,  -12'd123,  
12'd565,  12'd67,  12'd340,  -12'd29,  -12'd342,  12'd314,  12'd137,  12'd214,  -12'd335,  -12'd110,  -12'd247,  -12'd34,  12'd65,  -12'd282,  -12'd56,  12'd280,  
12'd340,  12'd223,  12'd248,  12'd146,  12'd110,  12'd213,  -12'd175,  12'd426,  -12'd258,  12'd132,  12'd39,  -12'd193,  12'd178,  12'd381,  12'd189,  -12'd20,  
-12'd197,  12'd29,  12'd447,  12'd97,  12'd24,  12'd108,  -12'd24,  12'd74,  12'd84,  12'd192,  -12'd199,  12'd141,  12'd45,  12'd299,  -12'd55,  -12'd269,  
-12'd348,  -12'd328,  -12'd32,  12'd40,  -12'd258,  -12'd92,  12'd317,  -12'd7,  -12'd261,  -12'd334,  -12'd105,  12'd88,  12'd24,  -12'd67,  12'd264,  12'd54,  
-12'd50,  12'd99,  -12'd8,  -12'd39,  12'd194,  -12'd372,  12'd126,  -12'd193,  -12'd100,  12'd501,  12'd169,  -12'd166,  -12'd159,  -12'd151,  -12'd179,  -12'd165,  
12'd190,  12'd109,  -12'd102,  12'd34,  12'd190,  -12'd175,  12'd82,  12'd396,  -12'd254,  -12'd258,  -12'd62,  12'd138,  -12'd186,  12'd225,  -12'd271,  12'd41,  

-12'd95,  12'd90,  -12'd269,  -12'd205,  12'd187,  12'd74,  12'd145,  -12'd29,  -12'd82,  12'd83,  12'd162,  12'd153,  -12'd54,  12'd318,  -12'd178,  -12'd141,  
12'd275,  -12'd125,  12'd18,  -12'd116,  -12'd231,  12'd13,  -12'd238,  -12'd73,  12'd243,  -12'd271,  -12'd194,  -12'd39,  -12'd0,  -12'd111,  -12'd331,  12'd2,  
12'd4,  -12'd76,  -12'd293,  -12'd73,  -12'd162,  12'd38,  -12'd378,  12'd35,  -12'd250,  12'd106,  -12'd239,  -12'd43,  12'd244,  -12'd443,  -12'd25,  12'd235,  
-12'd39,  12'd20,  -12'd251,  -12'd182,  -12'd134,  -12'd93,  12'd170,  -12'd118,  -12'd101,  -12'd401,  12'd77,  -12'd346,  12'd154,  -12'd281,  -12'd64,  -12'd198,  
-12'd444,  12'd89,  -12'd291,  12'd29,  12'd40,  12'd55,  12'd203,  12'd169,  12'd103,  12'd140,  -12'd89,  12'd94,  -12'd162,  -12'd347,  12'd229,  -12'd74,  
-12'd319,  -12'd194,  -12'd202,  -12'd226,  -12'd106,  12'd349,  12'd243,  -12'd8,  -12'd173,  12'd101,  -12'd13,  12'd18,  -12'd260,  12'd35,  -12'd311,  12'd217,  
12'd108,  -12'd349,  -12'd21,  -12'd109,  -12'd298,  -12'd157,  -12'd55,  12'd170,  -12'd8,  -12'd322,  -12'd236,  -12'd96,  -12'd127,  -12'd225,  12'd64,  12'd74,  
12'd124,  12'd269,  -12'd85,  -12'd125,  12'd279,  -12'd78,  -12'd36,  -12'd357,  12'd26,  -12'd30,  12'd56,  12'd39,  -12'd211,  -12'd26,  -12'd88,  -12'd112,  
-12'd114,  -12'd272,  -12'd408,  -12'd173,  -12'd300,  12'd327,  12'd53,  -12'd207,  12'd52,  12'd159,  -12'd2,  -12'd17,  -12'd458,  -12'd303,  -12'd278,  12'd169,  
12'd81,  -12'd212,  -12'd31,  -12'd269,  -12'd139,  12'd244,  -12'd38,  12'd50,  12'd167,  12'd251,  -12'd52,  -12'd13,  12'd136,  -12'd20,  -12'd66,  12'd201,  
-12'd65,  -12'd111,  12'd116,  12'd242,  12'd7,  -12'd215,  -12'd60,  -12'd16,  -12'd418,  12'd167,  -12'd60,  -12'd163,  -12'd78,  12'd69,  12'd163,  12'd73,  
-12'd202,  -12'd157,  -12'd73,  12'd85,  -12'd96,  12'd173,  12'd10,  -12'd397,  12'd52,  12'd123,  -12'd138,  12'd301,  -12'd135,  12'd236,  -12'd51,  12'd61,  
12'd41,  -12'd33,  12'd99,  -12'd63,  12'd2,  -12'd345,  -12'd98,  -12'd185,  -12'd57,  -12'd76,  -12'd62,  12'd56,  -12'd43,  -12'd267,  12'd25,  12'd215,  
12'd148,  -12'd207,  12'd55,  12'd147,  12'd208,  12'd28,  -12'd234,  -12'd99,  -12'd26,  -12'd150,  -12'd244,  -12'd32,  -12'd303,  12'd305,  12'd182,  -12'd123,  
12'd89,  -12'd24,  -12'd222,  -12'd248,  -12'd244,  -12'd207,  12'd99,  -12'd179,  12'd257,  -12'd192,  12'd161,  -12'd168,  12'd24,  12'd19,  12'd261,  12'd135,  
-12'd73,  -12'd103,  -12'd371,  12'd108,  -12'd43,  -12'd202,  -12'd434,  12'd111,  -12'd140,  12'd120,  -12'd367,  -12'd187,  -12'd173,  12'd142,  -12'd262,  -12'd75,  
-12'd140,  -12'd189,  12'd231,  12'd45,  -12'd113,  12'd57,  -12'd12,  -12'd78,  12'd46,  12'd72,  -12'd388,  12'd4,  -12'd227,  -12'd280,  12'd153,  -12'd239,  
-12'd156,  -12'd221,  -12'd269,  12'd116,  -12'd314,  12'd29,  -12'd93,  12'd211,  -12'd277,  -12'd140,  -12'd180,  12'd30,  -12'd265,  12'd78,  -12'd336,  12'd159,  
12'd156,  12'd71,  -12'd52,  12'd79,  -12'd5,  -12'd55,  12'd150,  -12'd139,  -12'd223,  -12'd119,  -12'd10,  -12'd111,  12'd170,  -12'd175,  -12'd207,  12'd28,  
12'd64,  12'd113,  -12'd50,  12'd173,  -12'd197,  -12'd2,  -12'd362,  -12'd28,  -12'd393,  12'd168,  -12'd225,  -12'd93,  12'd136,  -12'd153,  12'd373,  12'd327,  
12'd247,  -12'd175,  12'd71,  -12'd213,  -12'd172,  -12'd55,  12'd164,  -12'd200,  -12'd146,  -12'd180,  12'd257,  12'd287,  -12'd155,  -12'd325,  -12'd308,  12'd96,  
-12'd85,  12'd266,  -12'd158,  -12'd110,  -12'd95,  12'd44,  -12'd236,  -12'd10,  -12'd211,  12'd143,  -12'd38,  12'd5,  -12'd84,  -12'd393,  -12'd241,  -12'd367,  
12'd307,  -12'd19,  12'd277,  -12'd202,  -12'd98,  12'd94,  -12'd115,  -12'd237,  -12'd134,  -12'd12,  -12'd274,  -12'd146,  -12'd30,  12'd19,  -12'd13,  12'd48,  
-12'd208,  12'd101,  -12'd77,  12'd355,  -12'd372,  -12'd219,  -12'd95,  12'd108,  12'd223,  -12'd17,  -12'd155,  -12'd339,  12'd22,  -12'd267,  12'd277,  12'd129,  
12'd199,  12'd309,  12'd129,  12'd63,  -12'd191,  -12'd89,  -12'd141,  12'd69,  -12'd195,  -12'd1,  -12'd53,  -12'd168,  12'd233,  12'd138,  12'd224,  -12'd97,  

-12'd240,  -12'd347,  -12'd313,  -12'd111,  -12'd23,  -12'd115,  -12'd507,  12'd190,  12'd223,  12'd424,  12'd167,  -12'd26,  12'd289,  12'd149,  12'd207,  -12'd19,  
-12'd281,  12'd236,  12'd39,  12'd240,  -12'd130,  -12'd82,  -12'd338,  12'd293,  12'd12,  12'd245,  -12'd92,  -12'd5,  12'd145,  -12'd204,  12'd343,  -12'd193,  
-12'd167,  12'd160,  12'd285,  12'd416,  -12'd227,  12'd206,  -12'd17,  12'd118,  -12'd120,  -12'd357,  -12'd293,  12'd205,  12'd333,  -12'd525,  12'd321,  12'd205,  
-12'd104,  -12'd239,  12'd48,  12'd227,  12'd64,  -12'd154,  -12'd399,  12'd298,  -12'd165,  12'd370,  12'd82,  12'd59,  -12'd275,  -12'd712,  12'd548,  -12'd61,  
12'd219,  -12'd121,  12'd108,  12'd95,  -12'd77,  12'd201,  12'd142,  12'd221,  12'd299,  12'd323,  12'd130,  12'd34,  -12'd34,  -12'd82,  12'd110,  -12'd205,  
12'd120,  12'd345,  12'd290,  12'd78,  -12'd245,  12'd444,  -12'd14,  -12'd2,  12'd142,  -12'd255,  -12'd190,  12'd120,  12'd298,  -12'd21,  12'd36,  -12'd87,  
12'd307,  -12'd192,  12'd4,  -12'd80,  12'd11,  -12'd24,  -12'd155,  12'd155,  12'd198,  -12'd408,  -12'd104,  12'd231,  12'd149,  12'd358,  -12'd62,  12'd216,  
-12'd94,  12'd294,  12'd3,  -12'd308,  -12'd182,  12'd403,  12'd4,  -12'd81,  -12'd18,  -12'd157,  -12'd228,  -12'd150,  -12'd208,  12'd70,  12'd69,  12'd77,  
-12'd153,  12'd314,  12'd51,  -12'd74,  -12'd167,  12'd36,  -12'd238,  12'd87,  -12'd37,  12'd253,  -12'd32,  -12'd246,  -12'd127,  12'd253,  12'd178,  12'd262,  
-12'd236,  -12'd180,  -12'd178,  12'd91,  12'd134,  -12'd196,  12'd166,  -12'd190,  -12'd193,  12'd26,  -12'd22,  12'd89,  -12'd227,  -12'd316,  12'd172,  12'd241,  
12'd230,  -12'd63,  -12'd113,  12'd171,  12'd8,  12'd22,  -12'd194,  12'd269,  12'd366,  12'd152,  -12'd577,  -12'd67,  -12'd14,  12'd118,  12'd209,  -12'd26,  
12'd265,  -12'd108,  -12'd164,  -12'd333,  12'd128,  12'd214,  12'd244,  12'd52,  12'd165,  -12'd347,  -12'd203,  12'd44,  12'd408,  12'd97,  12'd227,  12'd270,  
-12'd239,  12'd432,  -12'd249,  -12'd362,  12'd130,  -12'd97,  12'd288,  -12'd76,  12'd99,  12'd230,  12'd112,  -12'd198,  12'd83,  12'd346,  -12'd70,  12'd100,  
12'd73,  12'd111,  12'd280,  12'd211,  -12'd18,  -12'd114,  -12'd24,  12'd72,  -12'd282,  -12'd179,  12'd50,  12'd82,  -12'd120,  12'd337,  12'd171,  12'd134,  
12'd46,  -12'd65,  12'd582,  -12'd194,  -12'd180,  12'd190,  12'd261,  -12'd292,  -12'd225,  -12'd175,  -12'd106,  12'd120,  -12'd390,  -12'd237,  12'd147,  12'd253,  
12'd68,  12'd80,  -12'd104,  12'd22,  12'd231,  12'd109,  12'd2,  -12'd171,  -12'd260,  12'd177,  -12'd529,  -12'd92,  12'd122,  12'd96,  -12'd45,  -12'd143,  
12'd60,  12'd178,  12'd119,  12'd89,  12'd343,  -12'd16,  12'd126,  12'd264,  -12'd13,  12'd97,  12'd278,  -12'd251,  12'd188,  -12'd245,  -12'd86,  12'd29,  
-12'd222,  12'd252,  -12'd99,  -12'd76,  -12'd221,  12'd133,  -12'd106,  -12'd132,  12'd188,  -12'd37,  -12'd235,  -12'd63,  -12'd89,  -12'd108,  -12'd83,  12'd83,  
12'd460,  12'd199,  12'd210,  12'd84,  12'd94,  12'd371,  -12'd16,  12'd14,  12'd267,  -12'd199,  12'd266,  12'd420,  12'd132,  -12'd225,  -12'd172,  -12'd69,  
12'd131,  12'd345,  -12'd79,  12'd13,  -12'd122,  -12'd53,  12'd126,  12'd97,  -12'd122,  -12'd15,  12'd20,  -12'd149,  12'd466,  -12'd116,  -12'd142,  12'd66,  
-12'd210,  12'd205,  -12'd144,  -12'd136,  -12'd75,  -12'd50,  -12'd251,  -12'd50,  -12'd23,  -12'd116,  -12'd123,  12'd231,  -12'd224,  -12'd135,  -12'd283,  -12'd53,  
-12'd9,  12'd34,  -12'd133,  12'd219,  12'd62,  12'd20,  12'd214,  -12'd172,  12'd5,  -12'd113,  12'd98,  12'd327,  -12'd251,  -12'd256,  -12'd112,  12'd381,  
-12'd361,  -12'd418,  12'd14,  -12'd289,  -12'd98,  -12'd38,  12'd165,  -12'd188,  -12'd309,  12'd183,  -12'd228,  12'd189,  12'd12,  -12'd155,  12'd54,  -12'd217,  
12'd340,  -12'd219,  12'd163,  -12'd119,  -12'd41,  -12'd187,  12'd169,  -12'd91,  -12'd121,  12'd188,  12'd66,  -12'd358,  12'd101,  12'd530,  -12'd470,  12'd194,  
-12'd246,  -12'd300,  -12'd82,  -12'd170,  12'd39,  -12'd135,  12'd171,  -12'd165,  -12'd107,  -12'd599,  -12'd474,  -12'd176,  12'd129,  -12'd167,  -12'd419,  12'd134,  

12'd162,  12'd116,  -12'd228,  12'd207,  12'd173,  12'd89,  12'd114,  -12'd93,  12'd69,  -12'd349,  12'd754,  12'd84,  -12'd141,  -12'd186,  -12'd187,  -12'd466,  
-12'd368,  -12'd275,  -12'd335,  12'd182,  -12'd315,  -12'd230,  -12'd523,  -12'd340,  12'd178,  -12'd145,  12'd279,  12'd108,  -12'd273,  -12'd201,  -12'd276,  -12'd228,  
12'd99,  12'd111,  -12'd109,  12'd218,  -12'd22,  12'd405,  -12'd442,  12'd369,  12'd73,  12'd62,  12'd31,  -12'd15,  -12'd221,  -12'd709,  -12'd215,  12'd342,  
-12'd432,  -12'd312,  12'd252,  -12'd331,  -12'd250,  12'd2,  -12'd22,  -12'd152,  12'd428,  12'd354,  12'd62,  -12'd170,  12'd201,  -12'd513,  -12'd32,  12'd72,  
-12'd108,  -12'd469,  12'd421,  -12'd54,  -12'd49,  -12'd353,  -12'd17,  12'd66,  12'd91,  12'd218,  12'd94,  -12'd203,  -12'd313,  -12'd90,  -12'd511,  12'd48,  
12'd264,  12'd11,  12'd136,  12'd334,  12'd80,  12'd258,  -12'd358,  12'd65,  12'd351,  12'd256,  12'd117,  12'd111,  12'd113,  -12'd40,  12'd24,  12'd34,  
12'd50,  12'd231,  12'd82,  -12'd104,  -12'd249,  12'd9,  -12'd170,  -12'd131,  12'd55,  -12'd32,  -12'd135,  -12'd106,  12'd44,  12'd11,  12'd106,  12'd303,  
12'd28,  -12'd174,  -12'd30,  12'd398,  -12'd190,  12'd91,  -12'd399,  12'd11,  -12'd81,  12'd161,  -12'd118,  12'd82,  -12'd220,  -12'd280,  12'd238,  12'd44,  
-12'd356,  12'd76,  -12'd203,  -12'd34,  -12'd171,  -12'd80,  12'd335,  -12'd172,  12'd252,  12'd276,  -12'd252,  -12'd351,  12'd83,  12'd43,  -12'd62,  -12'd113,  
-12'd325,  -12'd82,  -12'd233,  12'd268,  -12'd38,  -12'd63,  -12'd187,  12'd263,  -12'd27,  12'd291,  -12'd52,  -12'd92,  12'd32,  -12'd185,  -12'd429,  -12'd150,  
12'd88,  -12'd70,  -12'd7,  12'd127,  12'd333,  12'd120,  12'd54,  12'd282,  -12'd3,  12'd26,  12'd26,  -12'd158,  12'd152,  12'd98,  12'd218,  -12'd42,  
-12'd295,  12'd87,  -12'd5,  12'd362,  12'd290,  -12'd353,  -12'd79,  -12'd244,  12'd392,  -12'd174,  12'd440,  12'd2,  12'd138,  -12'd166,  12'd83,  12'd96,  
12'd140,  12'd226,  -12'd122,  12'd104,  -12'd51,  -12'd206,  -12'd7,  12'd264,  -12'd261,  -12'd30,  12'd312,  12'd115,  -12'd52,  -12'd256,  -12'd2,  12'd116,  
12'd421,  -12'd26,  12'd49,  -12'd252,  12'd73,  -12'd11,  12'd295,  12'd170,  -12'd166,  -12'd454,  12'd282,  -12'd74,  12'd71,  -12'd247,  12'd177,  12'd86,  
-12'd108,  12'd210,  12'd160,  -12'd68,  12'd297,  12'd331,  12'd153,  -12'd73,  -12'd67,  12'd188,  12'd120,  -12'd48,  12'd300,  12'd19,  -12'd197,  -12'd160,  
-12'd248,  12'd353,  12'd226,  12'd270,  12'd504,  -12'd160,  -12'd390,  12'd89,  -12'd12,  12'd59,  -12'd139,  -12'd134,  12'd153,  12'd4,  -12'd60,  12'd24,  
-12'd205,  12'd193,  -12'd104,  12'd227,  12'd298,  -12'd110,  -12'd504,  12'd134,  12'd317,  -12'd371,  12'd69,  -12'd114,  12'd160,  -12'd513,  12'd144,  -12'd5,  
12'd302,  -12'd302,  12'd288,  -12'd250,  -12'd262,  -12'd306,  -12'd168,  12'd8,  -12'd21,  -12'd18,  -12'd287,  12'd373,  -12'd142,  12'd454,  -12'd279,  -12'd125,  
12'd418,  12'd31,  12'd317,  -12'd209,  -12'd336,  -12'd109,  12'd340,  -12'd267,  12'd197,  -12'd86,  12'd95,  12'd356,  12'd208,  12'd74,  12'd82,  12'd128,  
-12'd92,  -12'd114,  -12'd475,  -12'd84,  -12'd94,  -12'd105,  -12'd192,  12'd323,  -12'd213,  12'd54,  12'd214,  12'd17,  -12'd98,  12'd32,  12'd298,  12'd267,  
-12'd343,  12'd482,  -12'd217,  -12'd355,  12'd75,  -12'd360,  12'd504,  -12'd269,  12'd261,  -12'd25,  -12'd259,  12'd60,  12'd125,  -12'd246,  -12'd62,  -12'd78,  
-12'd19,  -12'd87,  -12'd243,  -12'd169,  -12'd94,  12'd107,  12'd533,  12'd145,  12'd184,  -12'd376,  12'd131,  12'd100,  -12'd17,  -12'd230,  -12'd195,  -12'd291,  
-12'd341,  -12'd40,  -12'd62,  12'd42,  -12'd291,  -12'd242,  12'd245,  -12'd409,  12'd391,  12'd166,  12'd257,  -12'd25,  -12'd106,  12'd329,  12'd270,  12'd232,  
-12'd292,  -12'd190,  -12'd102,  12'd345,  12'd355,  -12'd238,  12'd245,  -12'd236,  -12'd44,  12'd84,  -12'd227,  12'd63,  -12'd57,  -12'd185,  12'd55,  -12'd74,  
-12'd252,  -12'd177,  12'd266,  -12'd33,  -12'd284,  12'd220,  12'd26,  -12'd91,  -12'd50,  12'd438,  -12'd281,  12'd267,  -12'd34,  12'd79,  12'd186,  12'd130,  

12'd163,  -12'd153,  12'd300,  -12'd250,  -12'd383,  -12'd193,  12'd98,  12'd0,  -12'd66,  12'd208,  12'd360,  -12'd169,  -12'd142,  -12'd32,  -12'd9,  -12'd174,  
-12'd306,  -12'd222,  -12'd532,  -12'd139,  -12'd86,  12'd73,  12'd148,  12'd176,  12'd265,  -12'd293,  12'd153,  12'd385,  12'd295,  -12'd329,  -12'd53,  -12'd41,  
12'd21,  12'd41,  -12'd381,  12'd200,  12'd434,  12'd256,  12'd22,  12'd120,  -12'd279,  12'd144,  12'd434,  12'd198,  12'd133,  -12'd209,  -12'd235,  -12'd145,  
12'd439,  12'd359,  12'd143,  12'd355,  -12'd30,  12'd176,  -12'd48,  12'd17,  12'd160,  12'd219,  12'd101,  -12'd23,  -12'd113,  -12'd549,  12'd13,  12'd216,  
-12'd16,  12'd143,  12'd6,  -12'd121,  12'd203,  12'd231,  12'd199,  12'd402,  -12'd153,  -12'd90,  12'd45,  -12'd173,  12'd506,  -12'd163,  -12'd329,  -12'd252,  
-12'd196,  -12'd379,  12'd158,  -12'd236,  12'd72,  -12'd36,  -12'd338,  -12'd95,  12'd388,  12'd166,  12'd208,  12'd237,  12'd22,  -12'd239,  12'd241,  -12'd372,  
12'd253,  12'd195,  12'd139,  -12'd367,  -12'd18,  -12'd377,  12'd153,  -12'd396,  -12'd311,  -12'd155,  12'd48,  -12'd65,  12'd130,  -12'd186,  -12'd198,  12'd70,  
-12'd215,  12'd32,  12'd146,  12'd213,  12'd257,  12'd210,  12'd413,  -12'd201,  -12'd326,  12'd49,  12'd242,  12'd229,  -12'd39,  -12'd368,  12'd352,  -12'd232,  
12'd210,  12'd95,  -12'd475,  12'd104,  12'd450,  12'd57,  12'd66,  12'd16,  12'd40,  -12'd180,  12'd237,  -12'd234,  12'd199,  -12'd225,  12'd266,  12'd110,  
-12'd800,  -12'd54,  -12'd505,  12'd181,  -12'd127,  -12'd264,  12'd12,  -12'd214,  12'd267,  12'd396,  12'd238,  12'd65,  12'd316,  12'd171,  -12'd11,  12'd444,  
12'd179,  -12'd41,  12'd121,  12'd262,  -12'd99,  -12'd28,  12'd321,  -12'd264,  -12'd246,  -12'd119,  -12'd374,  -12'd77,  -12'd92,  12'd90,  12'd322,  12'd241,  
12'd336,  -12'd135,  12'd123,  12'd293,  -12'd388,  12'd82,  12'd147,  -12'd82,  -12'd80,  -12'd404,  12'd450,  12'd80,  12'd144,  -12'd264,  12'd37,  -12'd288,  
12'd74,  -12'd357,  -12'd94,  12'd30,  -12'd135,  -12'd14,  12'd355,  12'd174,  12'd289,  12'd105,  12'd471,  -12'd243,  12'd318,  -12'd248,  12'd18,  -12'd50,  
12'd53,  12'd11,  -12'd126,  12'd106,  -12'd330,  12'd28,  -12'd257,  -12'd119,  12'd250,  -12'd278,  12'd130,  12'd63,  12'd45,  -12'd11,  12'd277,  12'd42,  
-12'd548,  -12'd246,  -12'd45,  12'd363,  -12'd103,  12'd75,  -12'd43,  -12'd59,  12'd101,  12'd767,  12'd385,  12'd300,  -12'd340,  12'd354,  -12'd36,  -12'd497,  
12'd14,  12'd141,  -12'd0,  12'd366,  -12'd54,  12'd130,  -12'd119,  -12'd68,  12'd185,  12'd260,  12'd231,  12'd324,  -12'd19,  -12'd238,  -12'd304,  12'd416,  
12'd418,  -12'd312,  12'd160,  12'd390,  -12'd115,  12'd170,  12'd633,  12'd371,  -12'd65,  -12'd408,  12'd128,  12'd26,  12'd348,  -12'd126,  12'd16,  12'd221,  
-12'd237,  12'd283,  -12'd71,  -12'd189,  -12'd117,  12'd103,  12'd142,  -12'd18,  12'd71,  -12'd45,  -12'd251,  12'd190,  -12'd140,  -12'd124,  -12'd107,  -12'd112,  
12'd294,  12'd42,  12'd345,  -12'd225,  -12'd510,  -12'd117,  12'd117,  12'd417,  12'd349,  12'd66,  12'd66,  -12'd144,  -12'd119,  -12'd102,  12'd39,  12'd214,  
12'd303,  -12'd88,  -12'd492,  12'd234,  12'd38,  -12'd343,  12'd82,  12'd254,  12'd398,  12'd104,  12'd113,  12'd148,  -12'd261,  12'd285,  12'd99,  -12'd78,  
12'd301,  12'd172,  -12'd18,  -12'd617,  -12'd253,  12'd116,  12'd180,  -12'd17,  -12'd525,  -12'd82,  12'd205,  12'd183,  -12'd260,  12'd17,  -12'd343,  12'd113,  
12'd158,  -12'd106,  12'd647,  -12'd68,  -12'd28,  -12'd68,  12'd422,  -12'd326,  12'd137,  12'd70,  -12'd207,  -12'd340,  12'd65,  12'd65,  -12'd219,  12'd335,  
-12'd100,  12'd170,  12'd62,  -12'd382,  12'd441,  -12'd127,  12'd257,  12'd41,  12'd597,  -12'd42,  -12'd319,  -12'd525,  -12'd301,  12'd581,  12'd266,  -12'd316,  
-12'd54,  -12'd501,  12'd111,  12'd81,  -12'd113,  -12'd312,  -12'd283,  -12'd446,  12'd494,  -12'd2,  -12'd358,  -12'd393,  -12'd547,  -12'd79,  -12'd42,  -12'd285,  
-12'd122,  -12'd440,  12'd6,  12'd14,  -12'd24,  12'd557,  12'd8,  -12'd92,  12'd197,  12'd489,  -12'd236,  -12'd152,  -12'd148,  12'd100,  12'd232,  -12'd33,  

12'd58,  -12'd370,  -12'd36,  -12'd45,  -12'd56,  12'd87,  -12'd135,  12'd337,  12'd443,  -12'd81,  -12'd84,  12'd124,  12'd153,  12'd99,  -12'd293,  -12'd60,  
12'd96,  12'd155,  12'd111,  -12'd336,  12'd173,  -12'd7,  12'd23,  12'd290,  12'd323,  -12'd26,  12'd276,  -12'd35,  -12'd8,  -12'd351,  12'd147,  -12'd216,  
12'd4,  -12'd146,  -12'd62,  12'd125,  12'd67,  12'd164,  -12'd200,  12'd5,  -12'd235,  12'd63,  -12'd101,  -12'd3,  -12'd39,  -12'd88,  12'd24,  -12'd101,  
-12'd32,  -12'd91,  -12'd79,  -12'd93,  -12'd36,  -12'd288,  12'd154,  12'd153,  12'd73,  -12'd11,  -12'd28,  -12'd6,  -12'd310,  -12'd39,  -12'd156,  -12'd68,  
-12'd89,  -12'd312,  12'd357,  -12'd151,  -12'd114,  -12'd11,  -12'd364,  -12'd30,  12'd234,  12'd68,  -12'd94,  12'd130,  -12'd29,  -12'd336,  12'd121,  -12'd19,  
-12'd167,  12'd236,  12'd107,  12'd53,  12'd8,  12'd199,  -12'd217,  -12'd19,  12'd234,  -12'd136,  -12'd145,  -12'd15,  12'd163,  -12'd364,  12'd278,  12'd35,  
-12'd86,  12'd55,  12'd0,  -12'd4,  -12'd101,  12'd215,  12'd186,  12'd120,  -12'd81,  -12'd238,  -12'd77,  -12'd194,  -12'd213,  12'd2,  -12'd292,  12'd283,  
12'd25,  -12'd189,  12'd309,  12'd216,  12'd107,  -12'd26,  -12'd351,  -12'd69,  -12'd341,  -12'd61,  -12'd79,  -12'd255,  12'd73,  -12'd224,  12'd166,  -12'd136,  
-12'd206,  -12'd214,  -12'd361,  12'd80,  -12'd40,  12'd4,  -12'd287,  12'd105,  -12'd33,  -12'd330,  12'd15,  -12'd48,  -12'd200,  -12'd73,  -12'd286,  -12'd265,  
-12'd26,  -12'd162,  12'd201,  12'd55,  12'd96,  -12'd84,  12'd0,  -12'd3,  -12'd351,  -12'd336,  12'd248,  -12'd101,  -12'd80,  12'd348,  12'd47,  -12'd158,  
-12'd9,  12'd20,  -12'd324,  -12'd80,  12'd153,  12'd122,  12'd116,  12'd97,  -12'd142,  12'd328,  12'd137,  -12'd235,  12'd95,  -12'd179,  -12'd52,  -12'd125,  
-12'd225,  12'd332,  -12'd219,  12'd200,  -12'd232,  12'd3,  -12'd124,  12'd66,  12'd64,  -12'd225,  -12'd187,  12'd175,  -12'd167,  12'd124,  -12'd437,  -12'd111,  
-12'd184,  -12'd28,  12'd35,  12'd201,  -12'd70,  12'd383,  -12'd301,  -12'd177,  -12'd216,  -12'd165,  -12'd4,  12'd135,  12'd48,  -12'd143,  12'd209,  -12'd241,  
12'd5,  12'd103,  -12'd244,  -12'd105,  12'd161,  -12'd165,  -12'd4,  -12'd298,  -12'd334,  -12'd297,  -12'd233,  -12'd327,  -12'd88,  12'd29,  12'd65,  -12'd164,  
12'd222,  12'd60,  12'd263,  12'd358,  -12'd293,  -12'd18,  12'd186,  -12'd145,  -12'd61,  12'd67,  -12'd109,  -12'd141,  12'd132,  -12'd61,  12'd81,  -12'd363,  
12'd237,  12'd92,  12'd84,  -12'd211,  12'd106,  12'd229,  12'd7,  12'd1,  12'd150,  12'd173,  -12'd104,  -12'd106,  -12'd195,  -12'd235,  -12'd350,  12'd1,  
12'd3,  -12'd222,  12'd111,  12'd43,  12'd148,  -12'd404,  -12'd274,  12'd121,  12'd78,  -12'd3,  12'd149,  -12'd41,  -12'd79,  -12'd239,  -12'd82,  -12'd208,  
12'd12,  -12'd135,  12'd1,  -12'd153,  12'd39,  -12'd103,  -12'd224,  -12'd321,  -12'd195,  12'd170,  12'd145,  -12'd115,  12'd98,  12'd329,  12'd58,  -12'd230,  
12'd4,  12'd233,  -12'd152,  -12'd294,  -12'd356,  -12'd292,  -12'd207,  -12'd160,  12'd80,  -12'd99,  12'd16,  -12'd257,  -12'd133,  12'd100,  -12'd124,  12'd73,  
-12'd291,  -12'd79,  -12'd33,  -12'd264,  12'd224,  12'd135,  12'd73,  -12'd125,  -12'd259,  -12'd198,  -12'd247,  -12'd288,  -12'd303,  12'd203,  -12'd40,  -12'd92,  
-12'd290,  -12'd21,  -12'd244,  12'd51,  12'd21,  12'd88,  -12'd94,  12'd110,  12'd281,  -12'd53,  12'd260,  -12'd30,  12'd134,  -12'd397,  12'd104,  12'd293,  
-12'd223,  -12'd179,  12'd336,  12'd98,  12'd8,  12'd297,  -12'd306,  -12'd98,  -12'd71,  12'd241,  -12'd203,  12'd147,  -12'd18,  -12'd85,  12'd42,  -12'd90,  
12'd73,  -12'd217,  -12'd121,  -12'd392,  12'd135,  -12'd202,  12'd147,  12'd4,  -12'd147,  12'd57,  -12'd109,  -12'd82,  12'd40,  -12'd161,  12'd47,  12'd17,  
-12'd176,  -12'd185,  12'd119,  12'd177,  -12'd270,  -12'd190,  -12'd65,  -12'd292,  -12'd132,  12'd46,  -12'd329,  -12'd328,  12'd29,  -12'd65,  -12'd60,  -12'd22,  
-12'd79,  12'd338,  12'd280,  -12'd48,  -12'd345,  12'd18,  -12'd51,  -12'd172,  -12'd142,  -12'd1,  -12'd412,  12'd222,  -12'd208,  -12'd204,  -12'd323,  -12'd13,  

-12'd196,  12'd25,  12'd417,  12'd400,  12'd12,  -12'd55,  -12'd255,  12'd358,  -12'd51,  12'd216,  12'd30,  -12'd552,  12'd286,  12'd205,  -12'd54,  12'd39,  
-12'd327,  -12'd11,  12'd454,  12'd196,  -12'd71,  -12'd228,  12'd20,  12'd145,  12'd181,  -12'd2,  12'd64,  -12'd134,  12'd157,  12'd932,  12'd218,  -12'd82,  
-12'd172,  -12'd92,  12'd558,  12'd28,  -12'd509,  -12'd21,  12'd231,  -12'd16,  -12'd64,  12'd192,  -12'd144,  12'd176,  -12'd113,  12'd721,  12'd61,  -12'd235,  
12'd514,  12'd137,  12'd222,  -12'd12,  12'd46,  12'd260,  12'd146,  -12'd287,  12'd395,  -12'd13,  12'd260,  12'd387,  -12'd229,  -12'd111,  -12'd17,  -12'd479,  
12'd473,  12'd623,  -12'd454,  12'd278,  -12'd324,  12'd208,  12'd329,  12'd196,  12'd124,  -12'd210,  12'd343,  -12'd62,  12'd340,  -12'd416,  -12'd147,  12'd506,  
-12'd51,  12'd278,  -12'd107,  -12'd330,  12'd540,  -12'd284,  -12'd256,  -12'd163,  -12'd311,  -12'd287,  12'd219,  12'd139,  12'd194,  12'd305,  12'd201,  -12'd201,  
-12'd193,  -12'd56,  12'd422,  12'd142,  -12'd86,  12'd246,  12'd196,  -12'd365,  -12'd150,  -12'd43,  12'd28,  12'd78,  12'd33,  12'd498,  12'd7,  -12'd29,  
-12'd85,  -12'd169,  12'd420,  12'd250,  -12'd206,  12'd213,  -12'd9,  -12'd188,  12'd326,  -12'd270,  -12'd25,  -12'd245,  -12'd203,  12'd584,  -12'd139,  -12'd320,  
12'd70,  -12'd172,  -12'd76,  12'd214,  -12'd198,  -12'd18,  12'd87,  12'd70,  -12'd40,  -12'd232,  -12'd162,  12'd92,  12'd251,  12'd122,  -12'd179,  -12'd169,  
12'd349,  -12'd200,  -12'd589,  12'd161,  12'd82,  -12'd230,  -12'd104,  -12'd153,  12'd381,  12'd293,  12'd155,  -12'd212,  -12'd176,  -12'd375,  -12'd252,  12'd258,  
-12'd15,  -12'd269,  12'd31,  12'd168,  -12'd66,  -12'd316,  -12'd176,  12'd63,  -12'd237,  -12'd108,  12'd124,  12'd92,  -12'd125,  -12'd156,  12'd189,  -12'd63,  
-12'd128,  -12'd107,  -12'd147,  -12'd187,  -12'd13,  -12'd89,  -12'd23,  -12'd32,  -12'd271,  -12'd119,  -12'd193,  -12'd160,  -12'd273,  12'd452,  -12'd82,  12'd293,  
12'd96,  -12'd219,  12'd372,  -12'd297,  -12'd314,  12'd220,  -12'd39,  12'd81,  -12'd210,  12'd213,  -12'd388,  -12'd63,  -12'd121,  12'd226,  12'd35,  12'd64,  
12'd287,  12'd121,  12'd390,  12'd425,  -12'd316,  12'd346,  -12'd85,  -12'd159,  12'd199,  -12'd468,  12'd1,  12'd49,  -12'd254,  12'd235,  -12'd320,  -12'd3,  
-12'd155,  -12'd339,  12'd225,  12'd303,  -12'd177,  12'd64,  -12'd176,  -12'd132,  12'd220,  -12'd83,  -12'd142,  -12'd266,  -12'd482,  -12'd250,  12'd178,  12'd101,  
-12'd286,  12'd246,  -12'd302,  12'd284,  12'd297,  12'd99,  12'd382,  12'd360,  12'd331,  12'd84,  12'd227,  -12'd263,  12'd259,  -12'd352,  -12'd335,  -12'd46,  
-12'd213,  -12'd317,  12'd136,  12'd57,  -12'd470,  -12'd378,  12'd151,  12'd114,  12'd46,  12'd502,  12'd203,  -12'd120,  12'd79,  -12'd174,  -12'd140,  12'd14,  
12'd83,  -12'd50,  -12'd134,  12'd239,  -12'd20,  12'd86,  12'd54,  12'd6,  -12'd8,  12'd136,  12'd14,  12'd25,  12'd228,  12'd436,  12'd74,  -12'd341,  
-12'd398,  -12'd47,  12'd84,  12'd325,  -12'd169,  -12'd246,  12'd159,  12'd337,  -12'd63,  -12'd244,  12'd337,  -12'd139,  12'd99,  -12'd162,  -12'd275,  12'd332,  
12'd184,  -12'd76,  12'd190,  12'd35,  12'd430,  -12'd111,  12'd86,  12'd21,  -12'd116,  -12'd151,  -12'd111,  12'd258,  12'd227,  12'd112,  12'd62,  12'd9,  
12'd9,  12'd234,  12'd98,  -12'd342,  -12'd376,  -12'd8,  12'd40,  -12'd290,  -12'd157,  12'd100,  12'd14,  12'd97,  -12'd195,  -12'd213,  12'd45,  12'd375,  
12'd121,  12'd252,  12'd469,  -12'd430,  12'd103,  12'd32,  12'd395,  -12'd108,  -12'd17,  12'd72,  12'd97,  12'd113,  12'd255,  12'd346,  12'd177,  -12'd19,  
-12'd24,  12'd141,  12'd138,  12'd124,  -12'd325,  -12'd63,  12'd160,  -12'd348,  -12'd11,  12'd15,  -12'd400,  -12'd205,  12'd334,  12'd422,  -12'd62,  12'd20,  
-12'd508,  12'd271,  -12'd556,  -12'd95,  12'd115,  -12'd43,  12'd128,  -12'd201,  -12'd211,  -12'd25,  12'd311,  -12'd638,  12'd42,  -12'd279,  12'd183,  12'd170,  
-12'd396,  12'd42,  -12'd354,  12'd11,  12'd34,  -12'd47,  -12'd62,  12'd227,  -12'd410,  -12'd499,  12'd107,  -12'd512,  -12'd305,  12'd274,  -12'd95,  -12'd69,  

-12'd484,  -12'd258,  12'd57,  -12'd197,  12'd614,  12'd98,  -12'd304,  12'd443,  -12'd142,  -12'd70,  12'd133,  -12'd177,  12'd10,  -12'd487,  -12'd48,  12'd13,  
12'd22,  12'd396,  12'd209,  -12'd44,  12'd307,  12'd199,  -12'd42,  12'd331,  -12'd133,  12'd329,  -12'd342,  -12'd234,  12'd292,  -12'd164,  12'd105,  12'd280,  
-12'd273,  -12'd214,  12'd243,  12'd116,  -12'd275,  12'd168,  12'd24,  -12'd232,  -12'd449,  12'd47,  -12'd218,  -12'd72,  12'd121,  12'd130,  12'd238,  12'd161,  
-12'd170,  12'd344,  12'd306,  12'd85,  12'd28,  12'd166,  12'd80,  12'd79,  12'd290,  12'd113,  12'd279,  12'd153,  -12'd398,  12'd562,  -12'd444,  12'd14,  
12'd464,  12'd396,  -12'd181,  12'd173,  -12'd1,  12'd247,  12'd254,  -12'd295,  12'd404,  -12'd117,  12'd203,  12'd62,  -12'd124,  12'd233,  12'd172,  12'd374,  
-12'd402,  -12'd29,  -12'd598,  -12'd174,  -12'd166,  -12'd70,  12'd73,  12'd133,  -12'd169,  -12'd31,  12'd395,  -12'd323,  -12'd299,  -12'd417,  -12'd251,  12'd118,  
-12'd366,  -12'd215,  -12'd234,  -12'd164,  12'd497,  -12'd103,  -12'd291,  12'd86,  -12'd133,  12'd25,  12'd99,  -12'd163,  -12'd280,  -12'd278,  -12'd255,  -12'd24,  
12'd287,  -12'd205,  12'd337,  12'd103,  12'd218,  -12'd123,  12'd117,  -12'd9,  -12'd545,  12'd211,  -12'd64,  12'd318,  -12'd29,  -12'd32,  -12'd160,  12'd44,  
12'd362,  -12'd56,  12'd452,  12'd139,  12'd344,  -12'd56,  12'd263,  12'd142,  12'd126,  -12'd315,  12'd184,  -12'd102,  12'd114,  12'd303,  12'd154,  -12'd109,  
12'd360,  -12'd23,  -12'd4,  12'd190,  -12'd15,  -12'd7,  12'd342,  12'd72,  12'd180,  12'd136,  -12'd105,  -12'd299,  12'd142,  -12'd151,  -12'd160,  12'd129,  
-12'd381,  -12'd252,  -12'd467,  -12'd274,  12'd199,  -12'd289,  -12'd288,  12'd138,  12'd419,  -12'd222,  12'd559,  -12'd15,  -12'd285,  -12'd313,  12'd107,  -12'd295,  
12'd135,  12'd97,  -12'd86,  12'd131,  -12'd41,  12'd248,  -12'd246,  12'd252,  -12'd103,  12'd1,  12'd4,  -12'd69,  -12'd209,  12'd177,  12'd191,  12'd59,  
12'd461,  -12'd212,  -12'd18,  -12'd331,  12'd67,  -12'd5,  -12'd261,  12'd216,  12'd176,  12'd267,  -12'd80,  -12'd69,  12'd413,  -12'd390,  -12'd212,  12'd93,  
12'd12,  -12'd355,  -12'd70,  12'd299,  12'd242,  -12'd91,  -12'd58,  12'd309,  -12'd209,  12'd334,  12'd145,  -12'd116,  12'd376,  -12'd16,  -12'd290,  12'd162,  
-12'd448,  12'd76,  -12'd189,  12'd177,  12'd145,  -12'd310,  12'd239,  -12'd244,  -12'd250,  12'd166,  12'd114,  12'd98,  -12'd2,  -12'd271,  12'd191,  12'd169,  
12'd167,  12'd112,  -12'd291,  12'd213,  -12'd273,  -12'd56,  -12'd78,  -12'd183,  12'd237,  -12'd203,  12'd93,  -12'd55,  -12'd195,  12'd328,  -12'd17,  -12'd219,  
12'd52,  -12'd198,  -12'd23,  12'd226,  -12'd278,  12'd126,  12'd48,  12'd58,  12'd169,  12'd196,  -12'd136,  -12'd239,  12'd201,  12'd373,  12'd383,  -12'd284,  
-12'd142,  12'd41,  12'd42,  12'd169,  12'd247,  12'd35,  12'd66,  -12'd180,  -12'd92,  -12'd260,  12'd319,  12'd313,  -12'd81,  12'd63,  -12'd200,  12'd258,  
-12'd64,  -12'd12,  -12'd143,  12'd141,  12'd46,  12'd170,  12'd218,  12'd77,  12'd261,  12'd300,  12'd159,  -12'd10,  -12'd315,  -12'd210,  12'd299,  12'd187,  
12'd114,  -12'd474,  -12'd340,  12'd64,  12'd258,  -12'd132,  -12'd202,  12'd110,  -12'd168,  12'd188,  12'd552,  12'd251,  12'd113,  12'd9,  -12'd149,  12'd379,  
12'd167,  -12'd34,  12'd365,  12'd361,  -12'd94,  -12'd43,  -12'd75,  -12'd104,  12'd218,  12'd20,  -12'd53,  -12'd13,  12'd91,  -12'd79,  12'd111,  12'd224,  
-12'd266,  -12'd142,  -12'd39,  12'd437,  12'd27,  12'd293,  -12'd262,  -12'd168,  -12'd298,  12'd253,  -12'd81,  -12'd61,  12'd81,  12'd298,  12'd305,  12'd108,  
12'd148,  12'd140,  12'd86,  -12'd21,  12'd69,  -12'd203,  -12'd257,  -12'd120,  -12'd252,  -12'd218,  -12'd52,  -12'd88,  12'd349,  -12'd133,  12'd155,  12'd324,  
-12'd26,  12'd283,  12'd112,  -12'd71,  -12'd177,  12'd13,  -12'd153,  -12'd211,  -12'd222,  -12'd302,  12'd295,  12'd24,  12'd184,  12'd123,  -12'd76,  12'd37,  
-12'd37,  12'd511,  12'd124,  -12'd228,  12'd258,  12'd21,  -12'd186,  12'd243,  -12'd205,  -12'd111,  12'd7,  -12'd57,  -12'd112,  12'd221,  -12'd51,  12'd90,  

-12'd137,  -12'd257,  -12'd293,  -12'd176,  12'd316,  12'd79,  12'd118,  12'd261,  -12'd244,  12'd210,  12'd275,  -12'd41,  12'd690,  -12'd99,  -12'd40,  -12'd294,  
12'd247,  -12'd95,  12'd8,  12'd216,  12'd41,  12'd217,  -12'd53,  12'd256,  -12'd228,  -12'd31,  12'd254,  12'd204,  12'd14,  12'd65,  12'd205,  12'd248,  
12'd487,  12'd133,  12'd125,  12'd185,  -12'd69,  12'd45,  -12'd152,  12'd122,  -12'd236,  -12'd358,  12'd177,  12'd11,  12'd138,  12'd101,  -12'd26,  12'd0,  
12'd34,  12'd126,  -12'd178,  12'd226,  -12'd60,  -12'd18,  -12'd1,  -12'd229,  -12'd257,  -12'd189,  12'd558,  -12'd17,  12'd366,  -12'd74,  -12'd89,  12'd25,  
-12'd44,  -12'd300,  -12'd346,  12'd391,  12'd231,  12'd115,  -12'd108,  12'd255,  -12'd62,  -12'd277,  12'd221,  -12'd244,  12'd252,  12'd297,  -12'd19,  -12'd166,  
12'd193,  12'd197,  -12'd265,  -12'd22,  12'd322,  -12'd132,  -12'd13,  -12'd63,  -12'd223,  -12'd186,  12'd345,  -12'd266,  12'd281,  -12'd216,  12'd11,  -12'd146,  
-12'd180,  12'd92,  -12'd186,  12'd117,  -12'd28,  12'd51,  12'd62,  12'd237,  -12'd206,  -12'd137,  12'd265,  -12'd399,  -12'd126,  -12'd269,  12'd9,  -12'd24,  
-12'd93,  12'd92,  12'd257,  12'd85,  12'd277,  12'd158,  -12'd72,  12'd172,  -12'd209,  12'd9,  12'd378,  -12'd199,  12'd222,  12'd650,  -12'd139,  12'd370,  
-12'd329,  12'd123,  12'd7,  -12'd12,  12'd27,  -12'd72,  -12'd38,  12'd282,  12'd317,  12'd145,  12'd401,  -12'd227,  -12'd48,  12'd60,  12'd205,  12'd137,  
12'd78,  12'd34,  12'd296,  -12'd57,  12'd97,  -12'd152,  12'd388,  12'd2,  12'd134,  -12'd70,  12'd458,  12'd360,  12'd44,  12'd123,  12'd56,  12'd87,  
-12'd321,  12'd452,  -12'd177,  -12'd241,  12'd151,  -12'd452,  -12'd96,  12'd70,  12'd411,  12'd77,  12'd595,  -12'd253,  12'd30,  12'd0,  -12'd66,  -12'd208,  
-12'd251,  -12'd135,  -12'd35,  -12'd232,  12'd205,  12'd67,  -12'd323,  -12'd15,  12'd75,  12'd418,  -12'd211,  -12'd91,  -12'd457,  -12'd313,  -12'd253,  -12'd42,  
12'd56,  -12'd52,  12'd102,  -12'd353,  12'd325,  12'd88,  -12'd96,  12'd17,  12'd180,  12'd430,  12'd123,  12'd347,  12'd186,  -12'd16,  12'd143,  12'd117,  
12'd188,  12'd65,  12'd134,  12'd98,  12'd223,  12'd161,  12'd59,  -12'd72,  12'd408,  -12'd97,  12'd70,  12'd356,  -12'd101,  12'd197,  12'd364,  12'd42,  
-12'd413,  12'd34,  -12'd425,  12'd66,  -12'd80,  -12'd580,  12'd20,  -12'd92,  12'd88,  12'd110,  -12'd14,  -12'd198,  12'd219,  12'd93,  12'd294,  -12'd156,  
12'd67,  -12'd336,  -12'd44,  -12'd24,  -12'd504,  12'd83,  -12'd55,  -12'd74,  12'd159,  -12'd314,  -12'd112,  -12'd94,  12'd74,  -12'd93,  -12'd230,  -12'd40,  
-12'd216,  -12'd347,  -12'd262,  12'd163,  -12'd436,  12'd108,  12'd159,  12'd192,  12'd245,  12'd292,  12'd108,  12'd408,  -12'd133,  12'd260,  12'd205,  -12'd324,  
-12'd104,  -12'd24,  12'd138,  12'd78,  12'd180,  12'd213,  12'd108,  -12'd12,  -12'd27,  -12'd144,  12'd269,  12'd71,  12'd228,  -12'd249,  12'd498,  -12'd380,  
-12'd283,  -12'd183,  12'd34,  12'd50,  12'd89,  12'd163,  12'd39,  -12'd9,  12'd107,  12'd38,  -12'd120,  -12'd40,  12'd73,  -12'd215,  -12'd20,  -12'd233,  
12'd33,  12'd153,  -12'd2,  -12'd105,  12'd127,  12'd46,  -12'd180,  12'd100,  -12'd87,  12'd230,  12'd26,  -12'd86,  -12'd330,  -12'd260,  -12'd253,  12'd197,  
-12'd84,  12'd86,  12'd62,  12'd93,  -12'd518,  12'd112,  -12'd9,  12'd26,  12'd534,  12'd111,  12'd107,  12'd98,  -12'd259,  12'd130,  12'd262,  -12'd74,  
12'd67,  -12'd272,  12'd5,  12'd215,  12'd141,  -12'd214,  -12'd37,  12'd210,  12'd204,  12'd156,  12'd287,  12'd144,  -12'd37,  12'd90,  -12'd29,  -12'd70,  
12'd312,  -12'd348,  -12'd254,  12'd152,  -12'd17,  12'd326,  12'd315,  12'd306,  12'd120,  12'd142,  -12'd179,  12'd43,  12'd227,  -12'd410,  12'd241,  12'd342,  
12'd25,  12'd364,  12'd103,  -12'd267,  12'd214,  -12'd93,  12'd56,  12'd12,  -12'd3,  12'd177,  12'd15,  -12'd97,  -12'd187,  12'd164,  -12'd145,  -12'd79,  
12'd269,  -12'd263,  12'd284,  12'd49,  -12'd391,  12'd237,  -12'd58,  12'd129,  12'd260,  12'd609,  -12'd138,  12'd146,  -12'd117,  12'd10,  -12'd221,  12'd290,  

12'd237,  -12'd353,  -12'd198,  -12'd122,  -12'd374,  12'd125,  12'd480,  -12'd354,  12'd249,  -12'd109,  -12'd49,  12'd285,  -12'd129,  -12'd22,  -12'd389,  -12'd404,  
-12'd235,  -12'd208,  -12'd474,  -12'd29,  -12'd0,  12'd161,  -12'd61,  -12'd170,  -12'd131,  12'd237,  -12'd218,  -12'd93,  -12'd289,  -12'd63,  12'd100,  -12'd34,  
-12'd278,  12'd60,  -12'd335,  -12'd152,  12'd454,  -12'd143,  -12'd442,  -12'd59,  -12'd32,  12'd70,  -12'd4,  -12'd169,  -12'd22,  -12'd887,  -12'd56,  12'd204,  
-12'd255,  -12'd207,  -12'd291,  -12'd16,  12'd141,  -12'd33,  -12'd370,  12'd163,  12'd162,  12'd205,  -12'd363,  12'd103,  -12'd194,  -12'd99,  -12'd215,  12'd92,  
-12'd371,  -12'd307,  12'd247,  12'd24,  -12'd16,  -12'd39,  -12'd197,  -12'd140,  -12'd70,  12'd230,  -12'd273,  -12'd146,  12'd352,  -12'd7,  12'd163,  12'd81,  
12'd9,  12'd120,  -12'd97,  -12'd120,  -12'd554,  12'd69,  12'd52,  12'd214,  12'd93,  12'd102,  12'd349,  -12'd23,  -12'd2,  -12'd115,  -12'd61,  12'd228,  
12'd182,  12'd172,  -12'd177,  -12'd164,  -12'd254,  12'd53,  12'd156,  -12'd100,  -12'd47,  12'd130,  -12'd266,  12'd144,  -12'd239,  12'd239,  12'd103,  12'd328,  
12'd229,  -12'd256,  -12'd410,  -12'd34,  12'd70,  12'd166,  12'd49,  -12'd43,  -12'd35,  12'd25,  -12'd189,  12'd35,  12'd320,  -12'd519,  12'd258,  -12'd38,  
-12'd5,  -12'd232,  -12'd413,  -12'd22,  12'd75,  -12'd222,  12'd171,  -12'd64,  12'd105,  -12'd215,  12'd116,  12'd27,  12'd156,  -12'd51,  -12'd73,  12'd162,  
-12'd436,  12'd61,  12'd379,  12'd20,  12'd22,  -12'd81,  12'd3,  12'd71,  -12'd275,  -12'd130,  12'd252,  -12'd265,  12'd110,  -12'd80,  12'd112,  -12'd117,  
-12'd122,  -12'd15,  12'd201,  12'd92,  12'd121,  -12'd64,  -12'd461,  12'd493,  12'd240,  -12'd72,  -12'd902,  -12'd223,  12'd226,  12'd351,  12'd303,  -12'd100,  
12'd56,  12'd165,  -12'd186,  12'd397,  12'd228,  12'd39,  -12'd272,  12'd166,  -12'd336,  -12'd172,  12'd209,  -12'd261,  12'd262,  12'd20,  12'd283,  -12'd147,  
12'd117,  12'd331,  -12'd434,  -12'd317,  12'd26,  12'd207,  12'd300,  -12'd148,  -12'd129,  -12'd164,  -12'd159,  12'd197,  -12'd31,  -12'd568,  -12'd221,  -12'd26,  
-12'd202,  12'd166,  12'd122,  -12'd594,  12'd232,  12'd99,  -12'd176,  12'd34,  -12'd79,  -12'd304,  -12'd45,  12'd76,  12'd8,  -12'd61,  -12'd254,  12'd322,  
12'd170,  12'd1,  12'd24,  -12'd250,  -12'd222,  12'd312,  -12'd106,  -12'd137,  12'd276,  12'd236,  12'd245,  -12'd68,  -12'd360,  12'd127,  -12'd4,  12'd175,  
-12'd32,  -12'd440,  -12'd135,  12'd436,  12'd327,  12'd257,  -12'd542,  12'd45,  -12'd117,  -12'd23,  -12'd171,  12'd16,  12'd243,  12'd61,  12'd1,  -12'd125,  
-12'd76,  -12'd154,  -12'd26,  -12'd30,  12'd569,  12'd76,  -12'd60,  -12'd122,  12'd30,  -12'd312,  12'd232,  -12'd65,  12'd287,  -12'd28,  -12'd42,  12'd3,  
12'd283,  12'd473,  12'd79,  -12'd48,  12'd456,  -12'd282,  12'd19,  12'd35,  -12'd336,  -12'd26,  12'd399,  -12'd238,  -12'd251,  12'd80,  -12'd237,  -12'd129,  
12'd160,  12'd276,  -12'd370,  -12'd138,  12'd394,  12'd310,  -12'd107,  -12'd106,  12'd318,  -12'd96,  -12'd254,  12'd329,  -12'd76,  12'd80,  -12'd236,  -12'd360,  
-12'd329,  -12'd515,  12'd99,  -12'd206,  -12'd325,  12'd54,  -12'd58,  12'd65,  12'd362,  -12'd3,  -12'd145,  -12'd369,  12'd257,  12'd174,  -12'd86,  -12'd352,  
12'd2,  12'd234,  -12'd84,  12'd317,  12'd426,  12'd192,  -12'd49,  12'd8,  12'd132,  12'd329,  12'd43,  12'd247,  12'd99,  -12'd369,  12'd449,  12'd44,  
12'd37,  -12'd126,  12'd99,  12'd263,  12'd245,  -12'd370,  12'd89,  -12'd41,  12'd257,  -12'd348,  12'd169,  12'd30,  12'd68,  -12'd224,  12'd12,  -12'd175,  
12'd309,  12'd18,  12'd200,  12'd257,  12'd42,  12'd306,  -12'd59,  -12'd127,  12'd434,  12'd157,  12'd237,  12'd300,  -12'd3,  -12'd306,  -12'd170,  12'd80,  
12'd251,  12'd162,  -12'd22,  -12'd107,  12'd78,  -12'd103,  -12'd113,  -12'd159,  12'd347,  -12'd126,  -12'd215,  12'd192,  12'd299,  12'd48,  12'd192,  -12'd166,  
12'd516,  -12'd259,  12'd370,  12'd136,  -12'd242,  12'd199,  12'd448,  -12'd146,  12'd717,  12'd161,  -12'd65,  12'd527,  12'd53,  12'd173,  12'd82,  -12'd211,  

-12'd221,  12'd209,  12'd278,  -12'd153,  12'd112,  12'd41,  12'd115,  12'd369,  12'd163,  -12'd131,  -12'd140,  12'd17,  12'd39,  12'd236,  -12'd270,  12'd483,  
-12'd68,  12'd263,  12'd475,  -12'd562,  12'd68,  -12'd231,  12'd370,  12'd115,  -12'd190,  -12'd16,  12'd2,  12'd152,  12'd75,  12'd258,  12'd32,  -12'd151,  
-12'd211,  12'd25,  12'd124,  -12'd185,  12'd237,  -12'd397,  12'd198,  -12'd223,  -12'd35,  -12'd146,  12'd297,  12'd400,  12'd341,  12'd770,  -12'd222,  12'd206,  
-12'd120,  12'd381,  12'd101,  -12'd160,  12'd319,  -12'd4,  12'd430,  12'd191,  -12'd28,  -12'd547,  -12'd121,  -12'd22,  12'd120,  12'd859,  -12'd155,  -12'd61,  
12'd237,  12'd102,  -12'd194,  -12'd70,  -12'd462,  12'd24,  12'd173,  -12'd142,  -12'd135,  -12'd163,  12'd57,  12'd126,  12'd284,  -12'd5,  -12'd142,  -12'd251,  
-12'd206,  -12'd65,  -12'd113,  12'd48,  12'd260,  -12'd210,  12'd26,  -12'd189,  -12'd266,  12'd219,  -12'd52,  -12'd242,  12'd35,  12'd384,  12'd143,  -12'd108,  
12'd302,  -12'd338,  12'd142,  12'd433,  -12'd149,  -12'd0,  12'd221,  -12'd12,  -12'd35,  -12'd190,  12'd267,  12'd126,  -12'd170,  12'd144,  -12'd237,  -12'd228,  
12'd365,  -12'd297,  12'd8,  12'd444,  -12'd18,  -12'd158,  12'd518,  -12'd194,  -12'd357,  -12'd30,  -12'd66,  12'd86,  -12'd143,  -12'd327,  -12'd339,  -12'd593,  
12'd505,  12'd354,  12'd325,  -12'd164,  -12'd8,  12'd69,  -12'd38,  -12'd29,  12'd332,  12'd228,  -12'd127,  12'd88,  12'd108,  12'd146,  -12'd125,  -12'd291,  
12'd577,  -12'd148,  -12'd160,  -12'd107,  12'd114,  -12'd38,  12'd252,  -12'd22,  12'd115,  12'd287,  -12'd39,  12'd263,  -12'd147,  -12'd47,  12'd36,  12'd91,  
-12'd175,  12'd49,  12'd225,  -12'd124,  12'd71,  12'd37,  12'd182,  12'd115,  -12'd19,  12'd64,  12'd152,  -12'd264,  -12'd150,  -12'd287,  -12'd218,  12'd385,  
12'd198,  12'd240,  -12'd65,  12'd355,  -12'd71,  -12'd157,  -12'd152,  12'd36,  -12'd167,  12'd162,  12'd156,  12'd104,  -12'd15,  12'd147,  12'd74,  -12'd60,  
-12'd36,  -12'd378,  -12'd175,  12'd54,  -12'd45,  12'd220,  -12'd190,  -12'd73,  -12'd55,  12'd55,  12'd70,  -12'd52,  -12'd24,  -12'd395,  -12'd87,  12'd252,  
-12'd95,  -12'd56,  12'd33,  12'd248,  12'd101,  12'd80,  -12'd5,  -12'd320,  12'd168,  12'd29,  -12'd0,  12'd318,  12'd29,  -12'd131,  -12'd18,  12'd397,  
-12'd181,  -12'd286,  12'd81,  12'd30,  12'd55,  12'd181,  -12'd143,  -12'd163,  12'd133,  12'd115,  12'd135,  12'd205,  -12'd81,  -12'd428,  12'd485,  12'd156,  
12'd114,  12'd301,  -12'd123,  -12'd119,  -12'd392,  -12'd90,  -12'd46,  -12'd30,  -12'd131,  -12'd83,  12'd198,  -12'd107,  12'd317,  -12'd25,  -12'd20,  12'd149,  
12'd30,  -12'd148,  12'd68,  12'd145,  12'd94,  12'd105,  -12'd98,  -12'd42,  -12'd62,  -12'd173,  -12'd423,  12'd250,  -12'd22,  -12'd118,  12'd118,  12'd42,  
12'd24,  12'd215,  -12'd123,  -12'd50,  12'd349,  12'd46,  -12'd172,  12'd266,  12'd62,  -12'd147,  12'd112,  12'd106,  -12'd208,  -12'd36,  -12'd185,  -12'd234,  
-12'd7,  -12'd95,  -12'd93,  12'd209,  -12'd106,  12'd142,  12'd298,  12'd48,  12'd60,  12'd1,  12'd163,  -12'd21,  12'd194,  -12'd166,  -12'd100,  12'd92,  
-12'd152,  12'd579,  -12'd25,  12'd138,  12'd229,  -12'd85,  12'd94,  -12'd7,  -12'd207,  -12'd285,  12'd98,  -12'd50,  -12'd21,  12'd325,  -12'd284,  12'd29,  
-12'd56,  12'd122,  12'd163,  -12'd567,  -12'd592,  12'd68,  12'd258,  -12'd166,  12'd157,  12'd92,  -12'd242,  -12'd256,  12'd50,  12'd406,  -12'd264,  -12'd142,  
-12'd125,  12'd167,  12'd197,  -12'd174,  -12'd18,  12'd240,  12'd218,  12'd28,  12'd10,  12'd197,  -12'd221,  12'd410,  -12'd117,  12'd323,  -12'd103,  12'd60,  
-12'd152,  12'd218,  12'd20,  -12'd187,  -12'd88,  12'd247,  12'd85,  12'd147,  12'd59,  -12'd321,  -12'd18,  -12'd39,  12'd175,  12'd40,  -12'd21,  -12'd428,  
-12'd110,  -12'd32,  -12'd314,  -12'd63,  12'd57,  -12'd114,  12'd210,  -12'd259,  12'd20,  -12'd47,  12'd15,  -12'd196,  -12'd33,  12'd216,  -12'd44,  12'd184,  
12'd406,  -12'd277,  -12'd306,  -12'd377,  -12'd338,  -12'd68,  12'd84,  -12'd88,  -12'd283,  -12'd596,  -12'd205,  -12'd669,  -12'd66,  -12'd95,  -12'd196,  -12'd412,  

-12'd36,  -12'd189,  12'd73,  12'd62,  -12'd108,  -12'd144,  12'd585,  -12'd189,  -12'd2,  -12'd22,  -12'd434,  12'd78,  -12'd556,  -12'd248,  12'd53,  -12'd7,  
-12'd421,  -12'd165,  12'd61,  -12'd276,  -12'd115,  -12'd111,  -12'd81,  -12'd478,  -12'd420,  -12'd74,  12'd253,  -12'd328,  -12'd161,  12'd14,  -12'd17,  -12'd154,  
-12'd131,  -12'd144,  12'd63,  -12'd311,  12'd75,  -12'd223,  12'd99,  12'd145,  12'd134,  12'd75,  12'd217,  -12'd127,  12'd89,  -12'd353,  12'd116,  12'd51,  
-12'd99,  12'd154,  12'd124,  12'd453,  -12'd126,  12'd285,  -12'd55,  12'd291,  12'd245,  -12'd30,  -12'd69,  12'd50,  -12'd90,  12'd64,  -12'd58,  -12'd217,  
12'd108,  12'd83,  -12'd78,  12'd541,  -12'd368,  12'd67,  -12'd197,  12'd80,  -12'd115,  -12'd10,  12'd52,  -12'd39,  12'd470,  12'd1,  12'd184,  -12'd50,  
-12'd63,  -12'd167,  -12'd127,  12'd175,  -12'd334,  -12'd166,  12'd283,  -12'd125,  12'd20,  12'd58,  12'd164,  -12'd301,  12'd40,  -12'd157,  12'd58,  -12'd23,  
12'd406,  -12'd289,  -12'd147,  12'd125,  -12'd163,  -12'd327,  -12'd25,  12'd122,  12'd244,  12'd47,  -12'd131,  -12'd17,  -12'd304,  12'd174,  12'd35,  -12'd337,  
-12'd17,  -12'd483,  -12'd122,  12'd78,  12'd292,  12'd42,  12'd43,  12'd78,  12'd454,  12'd301,  12'd264,  -12'd173,  12'd88,  -12'd4,  12'd382,  -12'd152,  
-12'd299,  12'd91,  -12'd133,  -12'd183,  12'd216,  -12'd273,  12'd37,  12'd446,  12'd182,  12'd8,  12'd160,  -12'd354,  12'd20,  -12'd508,  12'd38,  12'd216,  
-12'd474,  -12'd461,  12'd146,  -12'd98,  12'd193,  12'd22,  -12'd508,  12'd93,  12'd182,  12'd188,  -12'd0,  12'd17,  12'd396,  12'd94,  -12'd362,  -12'd15,  
-12'd71,  12'd114,  -12'd196,  12'd314,  12'd12,  12'd260,  -12'd23,  12'd286,  12'd82,  -12'd102,  -12'd635,  -12'd216,  12'd16,  12'd361,  12'd195,  12'd54,  
12'd6,  12'd65,  12'd140,  -12'd19,  -12'd337,  -12'd144,  -12'd240,  12'd227,  -12'd153,  12'd67,  -12'd81,  -12'd268,  -12'd165,  12'd167,  12'd100,  -12'd274,  
-12'd359,  -12'd24,  -12'd325,  -12'd5,  12'd176,  12'd154,  -12'd79,  -12'd78,  -12'd216,  12'd51,  12'd97,  -12'd402,  12'd133,  12'd9,  -12'd293,  12'd300,  
-12'd505,  -12'd179,  -12'd56,  -12'd158,  12'd220,  12'd260,  -12'd232,  12'd14,  12'd139,  12'd21,  12'd88,  -12'd240,  -12'd11,  -12'd343,  -12'd149,  12'd344,  
-12'd618,  -12'd140,  12'd381,  12'd218,  12'd189,  -12'd373,  12'd255,  -12'd279,  -12'd190,  12'd224,  -12'd229,  12'd151,  -12'd403,  12'd52,  12'd189,  -12'd67,  
-12'd112,  12'd178,  12'd66,  12'd427,  12'd95,  12'd353,  -12'd110,  -12'd3,  -12'd29,  12'd160,  -12'd28,  -12'd369,  12'd189,  12'd366,  -12'd78,  12'd226,  
-12'd198,  12'd218,  -12'd37,  12'd117,  12'd0,  12'd205,  -12'd196,  -12'd124,  -12'd222,  -12'd201,  12'd294,  -12'd27,  -12'd59,  12'd60,  12'd48,  -12'd39,  
12'd200,  12'd5,  -12'd197,  12'd67,  -12'd201,  -12'd287,  12'd181,  12'd249,  -12'd288,  12'd181,  12'd295,  12'd133,  12'd122,  12'd12,  -12'd114,  -12'd138,  
12'd81,  12'd449,  -12'd3,  -12'd435,  12'd37,  12'd158,  12'd145,  12'd175,  12'd309,  -12'd577,  -12'd10,  12'd223,  -12'd3,  12'd138,  -12'd153,  12'd119,  
12'd52,  12'd48,  12'd258,  -12'd239,  12'd156,  -12'd145,  12'd520,  12'd569,  -12'd19,  -12'd563,  -12'd202,  12'd19,  12'd79,  12'd147,  12'd125,  -12'd331,  
12'd168,  12'd185,  -12'd402,  12'd148,  12'd500,  12'd61,  12'd36,  12'd60,  12'd605,  12'd233,  12'd112,  12'd188,  -12'd242,  -12'd481,  -12'd203,  12'd209,  
-12'd43,  12'd105,  -12'd475,  12'd349,  -12'd13,  12'd210,  12'd70,  -12'd66,  12'd252,  12'd297,  12'd344,  12'd49,  -12'd180,  -12'd336,  -12'd173,  12'd98,  
12'd389,  12'd219,  12'd184,  12'd220,  12'd174,  -12'd112,  12'd84,  -12'd195,  12'd488,  -12'd47,  12'd138,  12'd303,  12'd99,  12'd190,  -12'd16,  12'd96,  
12'd258,  12'd6,  12'd196,  -12'd405,  -12'd56,  -12'd174,  12'd123,  12'd191,  12'd89,  12'd334,  -12'd25,  12'd428,  12'd212,  12'd450,  12'd90,  -12'd88,  
12'd270,  12'd16,  -12'd202,  -12'd277,  -12'd322,  12'd252,  12'd92,  -12'd179,  -12'd51,  -12'd186,  -12'd87,  12'd147,  12'd211,  12'd389,  -12'd45,  -12'd110,  

-12'd611,  12'd272,  12'd33,  -12'd363,  -12'd7,  12'd31,  12'd136,  -12'd424,  -12'd113,  -12'd428,  -12'd534,  12'd96,  -12'd485,  12'd162,  -12'd249,  12'd212,  
-12'd206,  12'd66,  12'd431,  12'd19,  12'd204,  -12'd246,  -12'd106,  -12'd241,  -12'd209,  -12'd241,  -12'd296,  12'd190,  -12'd178,  12'd31,  -12'd235,  -12'd41,  
12'd89,  12'd535,  -12'd80,  -12'd218,  12'd241,  12'd263,  -12'd264,  -12'd424,  12'd255,  12'd23,  -12'd89,  12'd129,  -12'd455,  12'd463,  -12'd38,  12'd108,  
12'd164,  12'd221,  -12'd152,  12'd31,  -12'd68,  12'd306,  -12'd14,  -12'd242,  12'd208,  -12'd75,  -12'd94,  -12'd191,  -12'd54,  12'd321,  -12'd165,  12'd200,  
12'd362,  12'd433,  -12'd464,  -12'd97,  12'd49,  12'd306,  12'd105,  -12'd147,  12'd28,  -12'd333,  12'd179,  12'd189,  12'd184,  -12'd160,  -12'd46,  -12'd76,  
12'd64,  12'd67,  12'd254,  -12'd58,  -12'd48,  -12'd11,  12'd201,  -12'd341,  -12'd580,  12'd157,  -12'd93,  12'd415,  -12'd329,  12'd223,  12'd287,  -12'd294,  
12'd55,  -12'd309,  12'd115,  -12'd125,  12'd175,  -12'd166,  12'd70,  -12'd10,  12'd256,  12'd1,  -12'd110,  12'd426,  -12'd144,  12'd137,  -12'd62,  -12'd323,  
12'd91,  12'd82,  12'd140,  -12'd137,  12'd195,  -12'd229,  12'd192,  -12'd232,  -12'd199,  12'd90,  -12'd120,  -12'd291,  12'd367,  -12'd137,  12'd344,  -12'd423,  
-12'd70,  -12'd406,  12'd144,  -12'd128,  12'd399,  -12'd100,  12'd60,  12'd162,  -12'd121,  -12'd183,  -12'd534,  12'd292,  -12'd373,  12'd19,  -12'd285,  12'd101,  
12'd131,  12'd264,  -12'd206,  -12'd304,  -12'd273,  -12'd124,  12'd230,  -12'd189,  12'd191,  -12'd139,  12'd355,  -12'd356,  -12'd34,  -12'd149,  -12'd29,  -12'd179,  
12'd51,  -12'd180,  12'd110,  12'd211,  -12'd375,  12'd42,  12'd59,  12'd139,  12'd143,  12'd222,  -12'd0,  -12'd122,  -12'd189,  12'd477,  12'd277,  -12'd225,  
-12'd10,  -12'd63,  12'd135,  12'd296,  -12'd201,  12'd385,  12'd80,  -12'd156,  12'd35,  12'd111,  -12'd300,  12'd148,  12'd252,  -12'd189,  -12'd64,  12'd134,  
12'd169,  -12'd95,  -12'd246,  12'd446,  12'd32,  -12'd45,  -12'd95,  12'd192,  -12'd290,  -12'd191,  12'd258,  -12'd235,  12'd246,  12'd147,  12'd357,  12'd220,  
12'd247,  -12'd163,  12'd517,  12'd99,  -12'd263,  12'd448,  12'd213,  12'd154,  12'd33,  -12'd330,  12'd23,  12'd66,  -12'd12,  -12'd131,  12'd58,  -12'd46,  
-12'd135,  -12'd142,  -12'd272,  12'd16,  -12'd37,  12'd64,  12'd33,  12'd70,  -12'd294,  -12'd171,  12'd77,  -12'd123,  12'd308,  12'd203,  -12'd88,  12'd159,  
12'd288,  -12'd209,  -12'd138,  12'd203,  12'd254,  12'd64,  12'd98,  12'd23,  -12'd298,  12'd155,  12'd215,  -12'd5,  12'd133,  12'd297,  12'd219,  12'd281,  
-12'd427,  12'd197,  12'd30,  12'd43,  12'd352,  -12'd271,  12'd192,  -12'd89,  12'd95,  12'd3,  12'd157,  12'd105,  12'd114,  -12'd78,  -12'd284,  12'd185,  
-12'd66,  12'd24,  -12'd124,  12'd171,  12'd7,  -12'd179,  -12'd56,  12'd69,  -12'd101,  -12'd11,  -12'd214,  -12'd292,  -12'd37,  -12'd224,  12'd178,  -12'd50,  
-12'd192,  12'd11,  -12'd157,  -12'd62,  -12'd11,  -12'd68,  -12'd94,  12'd417,  -12'd438,  -12'd184,  12'd143,  12'd145,  -12'd212,  -12'd333,  -12'd93,  -12'd187,  
12'd178,  -12'd221,  -12'd607,  -12'd8,  -12'd383,  12'd170,  -12'd131,  12'd90,  -12'd203,  -12'd211,  12'd51,  -12'd9,  -12'd84,  -12'd289,  12'd173,  12'd294,  
-12'd41,  12'd305,  12'd314,  12'd34,  12'd290,  12'd226,  -12'd68,  12'd286,  -12'd168,  -12'd274,  12'd165,  12'd239,  -12'd61,  -12'd211,  12'd25,  12'd19,  
12'd196,  12'd73,  12'd184,  -12'd81,  12'd332,  -12'd139,  12'd69,  -12'd235,  -12'd20,  -12'd52,  -12'd72,  -12'd89,  12'd2,  12'd156,  -12'd356,  12'd125,  
-12'd119,  12'd73,  -12'd188,  -12'd364,  12'd71,  -12'd315,  -12'd58,  -12'd150,  -12'd280,  12'd332,  -12'd129,  -12'd72,  -12'd61,  12'd336,  12'd101,  -12'd120,  
-12'd123,  12'd84,  12'd275,  12'd269,  12'd332,  -12'd260,  -12'd49,  -12'd55,  -12'd77,  12'd128,  12'd53,  12'd244,  12'd6,  12'd64,  -12'd117,  -12'd33,  
-12'd193,  -12'd284,  12'd119,  12'd422,  12'd113,  12'd106,  12'd158,  -12'd166,  -12'd290,  12'd398,  -12'd103,  12'd117,  -12'd128,  -12'd396,  12'd24,  12'd83,  

12'd4,  -12'd267,  -12'd72,  12'd150,  -12'd69,  -12'd39,  12'd40,  12'd142,  -12'd83,  -12'd41,  12'd604,  -12'd298,  12'd249,  -12'd141,  12'd69,  12'd363,  
12'd204,  -12'd13,  12'd100,  -12'd40,  -12'd173,  12'd322,  12'd44,  12'd48,  12'd17,  -12'd287,  12'd528,  -12'd10,  -12'd232,  -12'd311,  -12'd357,  -12'd168,  
-12'd94,  12'd163,  12'd187,  12'd105,  -12'd74,  -12'd147,  -12'd95,  -12'd165,  -12'd279,  -12'd306,  12'd304,  12'd138,  -12'd35,  -12'd57,  12'd3,  12'd395,  
12'd504,  -12'd94,  -12'd387,  -12'd96,  -12'd92,  -12'd211,  -12'd256,  12'd274,  12'd178,  12'd275,  12'd257,  -12'd52,  12'd9,  -12'd401,  -12'd20,  12'd45,  
12'd38,  12'd63,  12'd244,  12'd369,  -12'd82,  12'd204,  -12'd35,  12'd206,  12'd294,  12'd213,  12'd10,  -12'd69,  -12'd142,  12'd117,  12'd153,  12'd11,  
-12'd406,  12'd180,  12'd407,  12'd129,  12'd1,  -12'd298,  12'd44,  -12'd119,  -12'd143,  12'd136,  -12'd112,  12'd195,  -12'd527,  -12'd299,  12'd307,  12'd261,  
-12'd231,  12'd105,  -12'd140,  -12'd210,  -12'd83,  -12'd72,  12'd415,  -12'd284,  12'd123,  -12'd79,  12'd457,  -12'd67,  12'd72,  -12'd138,  -12'd536,  -12'd35,  
-12'd126,  12'd499,  12'd19,  12'd20,  12'd52,  12'd132,  12'd360,  -12'd299,  -12'd130,  -12'd58,  12'd197,  -12'd197,  12'd84,  12'd324,  -12'd512,  12'd0,  
-12'd182,  12'd244,  -12'd160,  -12'd129,  12'd261,  12'd141,  -12'd258,  12'd26,  12'd228,  -12'd21,  12'd399,  -12'd240,  12'd201,  12'd237,  12'd235,  12'd110,  
-12'd308,  -12'd334,  -12'd307,  12'd67,  12'd151,  -12'd101,  12'd154,  -12'd247,  12'd54,  -12'd64,  -12'd239,  -12'd70,  -12'd124,  12'd46,  12'd388,  -12'd29,  
12'd101,  -12'd214,  12'd159,  -12'd234,  -12'd296,  12'd311,  12'd45,  12'd152,  12'd100,  -12'd158,  -12'd435,  12'd109,  12'd2,  -12'd212,  12'd152,  -12'd117,  
12'd319,  -12'd20,  -12'd54,  12'd199,  12'd275,  12'd306,  -12'd146,  -12'd67,  12'd217,  12'd74,  12'd53,  -12'd52,  12'd40,  -12'd224,  12'd25,  -12'd10,  
12'd207,  -12'd89,  12'd32,  -12'd345,  -12'd145,  -12'd50,  -12'd219,  -12'd59,  12'd77,  12'd406,  -12'd203,  -12'd231,  12'd262,  12'd113,  -12'd378,  -12'd111,  
12'd282,  -12'd189,  -12'd22,  -12'd38,  12'd259,  12'd335,  12'd70,  -12'd262,  -12'd69,  -12'd256,  -12'd33,  12'd132,  -12'd774,  12'd295,  -12'd146,  12'd28,  
12'd97,  12'd132,  12'd659,  -12'd172,  -12'd404,  12'd20,  12'd409,  12'd176,  12'd253,  12'd301,  -12'd365,  12'd569,  -12'd350,  -12'd91,  -12'd241,  -12'd14,  
12'd312,  12'd318,  12'd325,  -12'd254,  -12'd316,  -12'd1,  -12'd87,  12'd313,  -12'd36,  -12'd97,  -12'd371,  12'd55,  -12'd87,  -12'd19,  -12'd78,  12'd47,  
-12'd89,  -12'd21,  12'd334,  12'd137,  -12'd277,  -12'd333,  12'd369,  -12'd126,  12'd132,  -12'd25,  12'd307,  12'd314,  12'd148,  12'd76,  -12'd69,  -12'd91,  
-12'd381,  -12'd178,  12'd306,  -12'd8,  -12'd248,  -12'd72,  12'd52,  -12'd26,  -12'd62,  12'd162,  12'd133,  12'd54,  -12'd110,  12'd306,  -12'd40,  12'd19,  
12'd450,  12'd292,  -12'd97,  12'd7,  -12'd339,  -12'd333,  12'd263,  12'd7,  12'd151,  12'd171,  12'd134,  12'd314,  12'd340,  12'd60,  -12'd94,  12'd50,  
12'd214,  12'd90,  12'd151,  12'd123,  12'd179,  12'd157,  -12'd162,  12'd277,  12'd319,  -12'd228,  12'd176,  12'd400,  12'd55,  12'd225,  12'd203,  12'd302,  
-12'd245,  12'd172,  12'd65,  -12'd250,  -12'd538,  12'd242,  12'd93,  12'd142,  -12'd520,  -12'd7,  -12'd120,  12'd251,  -12'd313,  12'd346,  -12'd324,  12'd218,  
12'd194,  12'd328,  -12'd246,  -12'd181,  -12'd39,  -12'd235,  12'd196,  -12'd63,  12'd365,  -12'd170,  -12'd178,  12'd5,  12'd161,  12'd265,  12'd410,  12'd121,  
-12'd203,  12'd58,  12'd219,  -12'd377,  -12'd203,  12'd65,  12'd141,  12'd130,  -12'd257,  -12'd111,  -12'd88,  -12'd218,  12'd203,  -12'd179,  12'd39,  12'd159,  
12'd38,  -12'd151,  12'd429,  -12'd111,  -12'd249,  -12'd394,  12'd284,  -12'd170,  -12'd134,  -12'd146,  12'd101,  -12'd49,  -12'd300,  12'd256,  -12'd20,  -12'd193,  
-12'd380,  -12'd161,  -12'd461,  -12'd346,  12'd18,  -12'd37,  -12'd147,  12'd69,  -12'd597,  -12'd293,  -12'd289,  -12'd539,  -12'd191,  12'd168,  -12'd326,  -12'd57,  

12'd41,  12'd93,  -12'd90,  12'd10,  12'd118,  12'd35,  -12'd6,  12'd384,  12'd46,  -12'd287,  12'd300,  -12'd22,  -12'd119,  -12'd109,  -12'd275,  -12'd171,  
12'd89,  12'd143,  12'd5,  12'd66,  12'd42,  12'd137,  12'd207,  12'd7,  -12'd246,  -12'd487,  -12'd375,  12'd90,  -12'd49,  12'd387,  12'd224,  12'd57,  
12'd302,  12'd149,  -12'd158,  12'd129,  -12'd203,  12'd49,  -12'd96,  -12'd324,  12'd389,  -12'd402,  -12'd148,  12'd223,  -12'd94,  12'd223,  -12'd47,  12'd39,  
-12'd117,  12'd88,  12'd199,  -12'd438,  12'd110,  -12'd47,  -12'd0,  12'd123,  12'd10,  12'd398,  12'd56,  -12'd5,  12'd225,  12'd384,  -12'd376,  12'd373,  
12'd48,  12'd167,  12'd88,  12'd102,  12'd79,  12'd115,  12'd259,  -12'd228,  12'd184,  12'd120,  12'd248,  12'd171,  12'd172,  -12'd350,  -12'd85,  12'd19,  
12'd35,  -12'd154,  -12'd491,  12'd263,  -12'd45,  -12'd28,  12'd76,  -12'd383,  -12'd1,  -12'd44,  -12'd185,  12'd39,  -12'd180,  -12'd170,  -12'd366,  -12'd91,  
12'd131,  12'd84,  12'd401,  12'd8,  -12'd309,  -12'd175,  -12'd363,  -12'd10,  -12'd129,  12'd15,  12'd219,  12'd209,  -12'd290,  12'd97,  12'd90,  12'd179,  
-12'd294,  -12'd358,  12'd161,  12'd224,  12'd65,  -12'd81,  -12'd168,  -12'd109,  -12'd118,  -12'd114,  12'd79,  -12'd117,  -12'd430,  -12'd25,  12'd330,  -12'd74,  
-12'd302,  12'd180,  -12'd58,  -12'd101,  -12'd11,  -12'd66,  -12'd84,  12'd21,  12'd86,  -12'd138,  -12'd264,  12'd119,  -12'd73,  12'd117,  12'd111,  -12'd120,  
12'd90,  12'd457,  12'd40,  12'd23,  -12'd49,  -12'd202,  -12'd93,  -12'd201,  12'd79,  12'd309,  -12'd370,  12'd316,  12'd78,  -12'd123,  -12'd154,  12'd238,  
12'd239,  12'd391,  -12'd303,  12'd57,  -12'd386,  12'd235,  -12'd97,  -12'd227,  12'd173,  -12'd219,  12'd324,  -12'd10,  -12'd18,  12'd36,  12'd351,  -12'd282,  
12'd112,  12'd251,  -12'd78,  12'd106,  -12'd71,  -12'd36,  -12'd76,  -12'd101,  12'd391,  12'd356,  12'd12,  12'd313,  12'd481,  12'd191,  -12'd392,  12'd27,  
-12'd58,  -12'd91,  -12'd9,  -12'd181,  -12'd155,  -12'd103,  12'd55,  12'd23,  12'd361,  -12'd33,  12'd44,  12'd208,  12'd190,  12'd2,  -12'd264,  -12'd135,  
-12'd169,  -12'd202,  12'd111,  12'd161,  -12'd210,  -12'd96,  -12'd172,  12'd30,  -12'd113,  12'd152,  -12'd273,  12'd136,  12'd152,  12'd279,  12'd34,  -12'd211,  
12'd436,  -12'd50,  -12'd482,  12'd110,  12'd81,  12'd475,  -12'd351,  -12'd65,  12'd329,  -12'd109,  12'd146,  -12'd61,  12'd118,  12'd165,  -12'd142,  12'd83,  
12'd384,  -12'd63,  12'd423,  12'd152,  -12'd192,  -12'd165,  12'd59,  -12'd153,  12'd41,  -12'd194,  -12'd208,  12'd26,  12'd208,  12'd239,  -12'd116,  12'd42,  
12'd406,  12'd270,  -12'd37,  12'd2,  -12'd147,  -12'd394,  -12'd16,  12'd27,  12'd269,  12'd46,  12'd56,  12'd423,  12'd309,  12'd118,  -12'd49,  12'd1,  
-12'd46,  12'd77,  -12'd137,  12'd47,  12'd109,  12'd231,  12'd60,  12'd168,  12'd215,  -12'd354,  12'd115,  -12'd127,  12'd217,  -12'd207,  -12'd214,  12'd143,  
-12'd102,  -12'd28,  -12'd26,  12'd358,  12'd523,  12'd247,  12'd149,  12'd96,  -12'd381,  12'd116,  -12'd81,  -12'd34,  -12'd259,  -12'd196,  12'd471,  12'd113,  
-12'd79,  -12'd241,  -12'd205,  12'd112,  -12'd212,  12'd66,  -12'd182,  12'd71,  -12'd88,  12'd524,  12'd356,  12'd328,  12'd228,  12'd284,  -12'd35,  12'd186,  
-12'd0,  -12'd248,  12'd357,  12'd92,  -12'd1,  12'd93,  12'd182,  12'd234,  -12'd186,  12'd34,  -12'd122,  -12'd386,  12'd14,  12'd366,  12'd315,  12'd32,  
-12'd118,  -12'd49,  -12'd254,  -12'd86,  -12'd52,  12'd66,  12'd228,  12'd126,  -12'd150,  -12'd357,  12'd43,  12'd118,  -12'd23,  -12'd155,  -12'd164,  -12'd175,  
-12'd246,  -12'd90,  12'd19,  12'd144,  12'd178,  -12'd163,  -12'd351,  -12'd12,  -12'd584,  -12'd268,  12'd227,  -12'd52,  -12'd185,  -12'd148,  -12'd218,  12'd74,  
-12'd483,  12'd58,  -12'd92,  12'd2,  -12'd7,  -12'd75,  -12'd95,  12'd130,  -12'd350,  12'd100,  -12'd186,  12'd52,  -12'd9,  -12'd195,  12'd32,  -12'd148,  
-12'd339,  -12'd50,  -12'd348,  12'd236,  12'd76,  -12'd119,  -12'd132,  12'd203,  12'd188,  12'd325,  12'd468,  12'd294,  12'd42,  12'd48,  12'd4,  12'd453,  

12'd175,  12'd218,  -12'd123,  -12'd229,  -12'd158,  -12'd122,  12'd52,  -12'd291,  -12'd240,  12'd0,  -12'd7,  12'd20,  -12'd264,  -12'd438,  -12'd316,  -12'd82,  
12'd307,  12'd120,  -12'd301,  12'd210,  -12'd264,  12'd113,  -12'd287,  12'd103,  12'd188,  -12'd94,  12'd198,  -12'd329,  -12'd40,  12'd19,  -12'd5,  -12'd17,  
12'd346,  -12'd171,  -12'd538,  12'd352,  -12'd182,  -12'd165,  -12'd146,  -12'd84,  12'd385,  12'd163,  -12'd303,  12'd106,  12'd168,  -12'd588,  -12'd62,  12'd513,  
-12'd109,  -12'd226,  12'd102,  -12'd106,  12'd316,  -12'd99,  -12'd435,  12'd46,  12'd6,  12'd324,  -12'd376,  -12'd53,  12'd61,  12'd112,  12'd192,  12'd193,  
-12'd28,  12'd12,  12'd249,  12'd83,  12'd238,  -12'd59,  -12'd418,  -12'd8,  -12'd190,  12'd239,  -12'd456,  -12'd108,  -12'd135,  12'd21,  -12'd227,  -12'd148,  
12'd115,  12'd28,  12'd129,  -12'd64,  12'd28,  12'd124,  -12'd152,  12'd63,  -12'd3,  12'd149,  -12'd115,  12'd244,  -12'd198,  12'd63,  -12'd143,  12'd105,  
-12'd73,  12'd257,  -12'd274,  -12'd113,  -12'd109,  -12'd172,  -12'd304,  12'd353,  -12'd114,  12'd139,  -12'd454,  12'd85,  12'd186,  12'd370,  12'd168,  12'd298,  
-12'd183,  -12'd306,  12'd140,  -12'd132,  12'd207,  12'd47,  -12'd179,  12'd102,  12'd36,  12'd250,  -12'd188,  12'd184,  -12'd55,  -12'd83,  12'd265,  -12'd136,  
-12'd70,  -12'd110,  12'd107,  12'd26,  -12'd254,  12'd96,  12'd78,  -12'd197,  -12'd290,  -12'd436,  -12'd125,  -12'd176,  12'd188,  12'd94,  12'd86,  -12'd128,  
12'd50,  -12'd114,  12'd38,  12'd270,  -12'd240,  -12'd79,  12'd88,  -12'd183,  12'd141,  -12'd532,  -12'd227,  -12'd102,  12'd169,  12'd75,  12'd65,  12'd50,  
12'd180,  12'd59,  -12'd219,  12'd92,  12'd438,  12'd176,  -12'd164,  -12'd92,  12'd211,  12'd424,  -12'd49,  12'd166,  12'd272,  12'd43,  12'd79,  -12'd195,  
-12'd204,  12'd157,  12'd297,  12'd94,  12'd49,  12'd309,  -12'd223,  12'd496,  -12'd203,  12'd177,  12'd85,  -12'd16,  12'd264,  12'd43,  12'd91,  -12'd64,  
12'd78,  12'd118,  12'd325,  -12'd1,  12'd127,  12'd29,  12'd428,  12'd159,  -12'd46,  -12'd192,  12'd2,  -12'd7,  12'd32,  12'd18,  12'd367,  -12'd299,  
12'd466,  12'd39,  12'd409,  -12'd44,  -12'd120,  12'd336,  12'd505,  -12'd117,  -12'd195,  -12'd24,  12'd269,  -12'd350,  -12'd197,  12'd303,  -12'd220,  -12'd58,  
12'd578,  12'd144,  -12'd506,  12'd85,  -12'd387,  12'd193,  12'd4,  12'd121,  -12'd50,  -12'd443,  -12'd319,  -12'd184,  12'd455,  12'd263,  -12'd69,  12'd303,  
-12'd418,  -12'd53,  -12'd335,  12'd99,  12'd782,  12'd292,  -12'd369,  -12'd168,  12'd38,  -12'd43,  -12'd157,  12'd158,  -12'd65,  -12'd324,  12'd183,  -12'd103,  
-12'd284,  12'd165,  12'd209,  12'd137,  12'd366,  -12'd111,  12'd25,  -12'd0,  -12'd26,  12'd150,  12'd230,  12'd48,  -12'd86,  12'd144,  -12'd470,  12'd140,  
12'd342,  -12'd201,  12'd236,  12'd88,  12'd81,  12'd217,  -12'd17,  12'd182,  12'd193,  -12'd64,  -12'd199,  12'd193,  -12'd69,  12'd97,  -12'd485,  -12'd97,  
-12'd126,  12'd171,  12'd218,  -12'd245,  -12'd33,  -12'd287,  12'd248,  -12'd164,  -12'd56,  12'd219,  -12'd289,  -12'd61,  -12'd297,  12'd276,  -12'd34,  12'd200,  
-12'd114,  -12'd201,  12'd52,  12'd276,  -12'd172,  -12'd126,  -12'd282,  -12'd81,  12'd61,  -12'd60,  -12'd385,  -12'd344,  -12'd180,  12'd451,  -12'd102,  -12'd164,  
-12'd92,  12'd27,  -12'd166,  12'd174,  12'd357,  -12'd179,  -12'd71,  -12'd147,  12'd225,  -12'd92,  12'd20,  -12'd82,  12'd92,  12'd10,  12'd121,  12'd66,  
-12'd166,  -12'd323,  -12'd0,  12'd309,  12'd89,  -12'd71,  12'd395,  12'd309,  12'd437,  12'd142,  12'd342,  -12'd239,  12'd11,  12'd59,  12'd55,  12'd198,  
-12'd223,  12'd40,  12'd23,  12'd152,  -12'd56,  -12'd20,  -12'd154,  -12'd310,  -12'd124,  -12'd73,  12'd5,  12'd24,  12'd43,  12'd189,  -12'd159,  12'd220,  
-12'd214,  -12'd343,  12'd92,  -12'd101,  12'd124,  -12'd21,  12'd147,  12'd224,  12'd151,  12'd75,  -12'd11,  -12'd284,  12'd37,  12'd200,  12'd226,  12'd258,  
-12'd88,  -12'd385,  12'd125,  -12'd11,  -12'd186,  12'd171,  -12'd13,  -12'd375,  12'd113,  -12'd108,  -12'd161,  12'd322,  12'd324,  12'd340,  12'd225,  12'd55,  

-12'd23,  12'd4,  -12'd300,  -12'd51,  -12'd3,  -12'd57,  -12'd101,  -12'd24,  -12'd341,  12'd87,  12'd189,  -12'd198,  -12'd34,  12'd190,  -12'd205,  12'd26,  
12'd62,  12'd42,  -12'd187,  12'd279,  -12'd125,  -12'd142,  12'd140,  -12'd261,  12'd306,  -12'd240,  12'd229,  -12'd350,  12'd240,  12'd61,  12'd139,  -12'd74,  
-12'd121,  12'd76,  -12'd161,  -12'd253,  -12'd120,  12'd180,  -12'd359,  -12'd220,  -12'd257,  12'd308,  -12'd303,  -12'd157,  12'd54,  -12'd36,  -12'd0,  -12'd75,  
-12'd152,  -12'd140,  -12'd97,  -12'd112,  -12'd50,  -12'd110,  -12'd182,  -12'd97,  -12'd162,  12'd212,  12'd226,  -12'd164,  -12'd43,  -12'd2,  12'd16,  12'd134,  
12'd7,  -12'd271,  -12'd12,  12'd172,  12'd213,  12'd128,  -12'd118,  12'd160,  12'd194,  12'd88,  12'd260,  -12'd147,  12'd182,  -12'd240,  -12'd24,  12'd186,  
12'd121,  -12'd45,  -12'd23,  12'd185,  -12'd205,  -12'd326,  -12'd117,  -12'd140,  12'd152,  12'd365,  12'd100,  12'd122,  12'd12,  -12'd34,  12'd319,  -12'd86,  
-12'd88,  -12'd35,  -12'd150,  -12'd125,  -12'd24,  -12'd373,  -12'd22,  12'd113,  -12'd15,  12'd85,  -12'd63,  -12'd151,  12'd144,  -12'd88,  -12'd158,  -12'd144,  
-12'd209,  12'd333,  -12'd50,  12'd64,  12'd214,  12'd67,  12'd72,  12'd33,  -12'd190,  12'd15,  -12'd38,  -12'd184,  -12'd136,  -12'd188,  -12'd50,  -12'd203,  
12'd277,  -12'd24,  12'd278,  12'd101,  12'd106,  -12'd283,  -12'd218,  -12'd43,  12'd136,  -12'd204,  -12'd52,  -12'd279,  12'd96,  12'd241,  -12'd114,  -12'd295,  
12'd117,  12'd180,  12'd21,  12'd242,  -12'd16,  -12'd138,  -12'd262,  -12'd189,  -12'd365,  12'd90,  -12'd247,  -12'd172,  -12'd206,  12'd156,  -12'd83,  12'd186,  
12'd268,  -12'd427,  12'd169,  -12'd338,  -12'd118,  12'd207,  12'd81,  -12'd242,  -12'd132,  12'd92,  -12'd49,  -12'd179,  12'd221,  -12'd133,  -12'd122,  -12'd187,  
12'd357,  -12'd8,  -12'd64,  -12'd100,  -12'd101,  -12'd135,  12'd241,  -12'd51,  -12'd83,  -12'd124,  -12'd177,  -12'd25,  12'd85,  12'd106,  12'd142,  -12'd404,  
12'd261,  12'd145,  12'd51,  -12'd378,  12'd65,  12'd64,  -12'd421,  12'd35,  12'd35,  12'd297,  12'd197,  -12'd32,  12'd32,  12'd19,  12'd9,  12'd193,  
-12'd129,  12'd291,  -12'd333,  -12'd1,  -12'd215,  -12'd37,  -12'd156,  12'd135,  -12'd119,  12'd131,  12'd261,  -12'd259,  -12'd72,  -12'd100,  -12'd15,  12'd178,  
-12'd191,  -12'd35,  -12'd267,  -12'd400,  -12'd150,  12'd215,  -12'd94,  -12'd81,  12'd129,  -12'd36,  12'd114,  -12'd148,  -12'd96,  12'd47,  -12'd140,  -12'd292,  
-12'd153,  12'd54,  12'd46,  -12'd226,  12'd96,  -12'd254,  12'd332,  12'd167,  -12'd270,  12'd74,  12'd22,  12'd187,  -12'd74,  12'd9,  -12'd44,  -12'd122,  
12'd317,  12'd136,  12'd56,  -12'd227,  -12'd168,  -12'd107,  12'd204,  -12'd300,  12'd183,  -12'd8,  -12'd110,  -12'd163,  -12'd121,  -12'd287,  12'd35,  -12'd226,  
-12'd111,  -12'd86,  -12'd254,  12'd341,  -12'd31,  12'd375,  -12'd123,  -12'd185,  -12'd322,  12'd24,  -12'd317,  -12'd192,  -12'd184,  -12'd136,  -12'd178,  -12'd179,  
-12'd98,  12'd121,  12'd123,  12'd10,  -12'd62,  -12'd335,  12'd31,  12'd288,  12'd90,  -12'd158,  -12'd56,  12'd6,  12'd87,  -12'd68,  12'd90,  12'd193,  
-12'd267,  -12'd159,  12'd259,  12'd63,  -12'd7,  -12'd77,  -12'd147,  -12'd143,  -12'd321,  12'd154,  12'd133,  12'd177,  12'd310,  -12'd27,  -12'd226,  12'd104,  
-12'd59,  -12'd228,  12'd222,  12'd272,  -12'd95,  -12'd17,  -12'd423,  12'd249,  -12'd170,  -12'd184,  -12'd308,  -12'd209,  -12'd31,  -12'd204,  -12'd159,  -12'd192,  
-12'd10,  -12'd259,  -12'd23,  12'd4,  -12'd330,  -12'd78,  -12'd335,  -12'd45,  -12'd15,  -12'd135,  12'd311,  -12'd137,  -12'd326,  12'd47,  -12'd138,  -12'd142,  
-12'd302,  -12'd129,  12'd9,  12'd26,  12'd21,  -12'd227,  -12'd23,  -12'd313,  -12'd246,  12'd118,  -12'd215,  12'd241,  12'd17,  -12'd146,  12'd289,  -12'd268,  
12'd40,  12'd16,  -12'd57,  12'd250,  -12'd92,  12'd103,  -12'd154,  12'd153,  -12'd103,  -12'd147,  -12'd72,  -12'd182,  12'd109,  -12'd404,  -12'd33,  -12'd346,  
12'd268,  -12'd138,  -12'd225,  -12'd347,  -12'd127,  12'd196,  -12'd67,  -12'd26,  -12'd118,  -12'd107,  12'd68,  12'd97,  12'd244,  -12'd269,  12'd177,  12'd146,  

-12'd69,  12'd46,  12'd252,  12'd74,  -12'd204,  -12'd187,  12'd162,  12'd313,  12'd70,  12'd59,  -12'd4,  -12'd106,  12'd219,  12'd268,  -12'd1,  12'd94,  
-12'd144,  12'd44,  12'd663,  -12'd498,  12'd284,  -12'd326,  12'd267,  12'd6,  -12'd182,  12'd33,  -12'd652,  12'd79,  -12'd2,  12'd515,  -12'd48,  12'd57,  
12'd116,  12'd78,  12'd0,  -12'd377,  12'd19,  -12'd242,  12'd575,  12'd85,  -12'd175,  12'd5,  -12'd207,  -12'd85,  -12'd322,  12'd677,  -12'd250,  -12'd367,  
-12'd221,  12'd190,  12'd183,  -12'd148,  12'd233,  -12'd118,  12'd354,  -12'd249,  12'd82,  -12'd90,  12'd59,  -12'd160,  -12'd375,  12'd350,  12'd274,  -12'd286,  
12'd291,  12'd253,  -12'd244,  -12'd93,  12'd8,  12'd550,  12'd114,  12'd64,  12'd191,  12'd88,  12'd58,  -12'd127,  12'd121,  -12'd110,  -12'd64,  12'd112,  
12'd9,  -12'd116,  12'd18,  12'd148,  12'd135,  12'd45,  12'd110,  -12'd46,  -12'd309,  -12'd154,  -12'd180,  12'd221,  12'd39,  12'd182,  12'd40,  -12'd156,  
12'd319,  -12'd353,  12'd111,  12'd129,  -12'd136,  -12'd364,  12'd273,  -12'd10,  -12'd51,  -12'd170,  -12'd260,  12'd149,  -12'd351,  12'd503,  -12'd297,  -12'd430,  
12'd19,  12'd255,  12'd294,  -12'd81,  -12'd236,  -12'd160,  12'd196,  -12'd152,  12'd150,  12'd20,  -12'd93,  -12'd49,  -12'd185,  12'd392,  12'd135,  -12'd478,  
12'd192,  -12'd47,  -12'd131,  -12'd413,  12'd275,  -12'd231,  -12'd89,  -12'd59,  -12'd113,  -12'd479,  -12'd117,  12'd128,  12'd120,  12'd174,  -12'd367,  -12'd31,  
12'd352,  12'd68,  12'd94,  -12'd239,  12'd26,  12'd286,  12'd85,  -12'd156,  12'd445,  12'd41,  12'd161,  -12'd113,  -12'd156,  -12'd55,  -12'd127,  -12'd162,  
-12'd179,  -12'd167,  -12'd453,  12'd102,  -12'd251,  12'd30,  12'd111,  -12'd200,  -12'd61,  -12'd156,  12'd497,  12'd111,  12'd357,  12'd158,  12'd109,  -12'd191,  
12'd91,  12'd35,  12'd32,  12'd68,  -12'd408,  12'd62,  12'd242,  -12'd246,  -12'd42,  12'd267,  -12'd109,  -12'd199,  12'd328,  12'd105,  12'd104,  12'd330,  
-12'd170,  12'd74,  12'd83,  12'd312,  12'd246,  12'd9,  12'd11,  -12'd36,  -12'd105,  -12'd154,  12'd268,  -12'd94,  12'd313,  -12'd160,  -12'd10,  -12'd95,  
-12'd159,  -12'd414,  12'd155,  12'd103,  12'd209,  12'd205,  12'd127,  12'd123,  12'd326,  -12'd234,  12'd21,  -12'd85,  -12'd136,  -12'd383,  -12'd37,  12'd138,  
-12'd214,  -12'd24,  -12'd265,  12'd252,  -12'd60,  12'd60,  -12'd33,  -12'd271,  -12'd330,  12'd252,  12'd53,  -12'd70,  12'd206,  -12'd258,  -12'd27,  12'd130,  
-12'd236,  12'd37,  12'd187,  -12'd276,  -12'd222,  -12'd147,  -12'd256,  -12'd9,  12'd181,  -12'd81,  12'd52,  12'd57,  12'd445,  -12'd9,  12'd210,  -12'd136,  
12'd58,  -12'd112,  -12'd20,  -12'd50,  12'd59,  12'd22,  12'd203,  12'd260,  -12'd151,  12'd107,  12'd343,  12'd336,  -12'd55,  12'd160,  -12'd143,  12'd82,  
12'd191,  -12'd314,  -12'd318,  12'd321,  12'd30,  12'd411,  -12'd91,  -12'd57,  -12'd329,  -12'd186,  12'd120,  12'd72,  12'd23,  12'd147,  12'd169,  -12'd40,  
-12'd8,  12'd25,  12'd206,  12'd351,  -12'd149,  12'd36,  12'd44,  12'd431,  12'd134,  12'd270,  12'd257,  12'd176,  -12'd183,  -12'd37,  12'd265,  12'd200,  
12'd5,  12'd93,  -12'd211,  12'd111,  12'd46,  -12'd209,  -12'd214,  -12'd148,  -12'd65,  -12'd162,  12'd262,  -12'd67,  12'd216,  12'd53,  12'd190,  12'd212,  
-12'd28,  -12'd126,  12'd175,  -12'd76,  -12'd163,  -12'd60,  -12'd30,  -12'd1,  -12'd254,  12'd166,  -12'd462,  -12'd248,  12'd79,  12'd38,  12'd237,  -12'd145,  
-12'd134,  12'd8,  12'd123,  -12'd106,  -12'd195,  -12'd208,  12'd189,  12'd36,  12'd65,  12'd96,  12'd51,  12'd82,  -12'd397,  12'd178,  -12'd115,  -12'd108,  
12'd302,  12'd474,  -12'd30,  -12'd49,  12'd220,  -12'd94,  -12'd182,  -12'd167,  -12'd532,  12'd42,  12'd33,  -12'd52,  -12'd390,  12'd170,  -12'd219,  -12'd185,  
-12'd290,  12'd421,  12'd276,  12'd248,  12'd372,  12'd19,  -12'd120,  -12'd57,  12'd277,  12'd489,  -12'd109,  -12'd281,  12'd19,  -12'd84,  12'd366,  -12'd126,  
12'd9,  -12'd115,  -12'd217,  12'd113,  12'd296,  12'd149,  12'd103,  12'd278,  -12'd63,  12'd371,  12'd194,  12'd49,  -12'd274,  12'd42,  12'd178,  12'd368,  

-12'd504,  -12'd8,  12'd39,  12'd74,  12'd90,  12'd153,  12'd21,  -12'd125,  12'd137,  12'd133,  12'd374,  -12'd354,  -12'd41,  -12'd114,  12'd552,  -12'd57,  
-12'd277,  -12'd290,  -12'd380,  -12'd133,  12'd132,  -12'd191,  -12'd225,  12'd291,  12'd173,  12'd25,  12'd142,  -12'd128,  12'd90,  12'd90,  12'd6,  12'd102,  
12'd53,  -12'd652,  12'd285,  12'd295,  12'd275,  -12'd274,  12'd27,  12'd175,  -12'd110,  -12'd59,  12'd97,  12'd246,  -12'd133,  -12'd306,  12'd255,  -12'd312,  
12'd55,  -12'd371,  12'd111,  12'd142,  -12'd233,  12'd204,  12'd165,  -12'd46,  12'd183,  -12'd63,  12'd140,  12'd103,  -12'd199,  -12'd13,  -12'd106,  -12'd183,  
-12'd421,  -12'd246,  12'd214,  -12'd130,  -12'd214,  12'd61,  -12'd80,  12'd282,  -12'd186,  12'd228,  -12'd203,  -12'd184,  -12'd45,  -12'd60,  -12'd91,  -12'd326,  
12'd72,  12'd180,  12'd71,  -12'd218,  -12'd175,  -12'd179,  -12'd437,  12'd142,  -12'd331,  12'd142,  12'd79,  12'd283,  -12'd229,  12'd211,  -12'd290,  -12'd381,  
-12'd190,  -12'd176,  -12'd466,  -12'd232,  12'd191,  12'd151,  12'd170,  -12'd457,  -12'd174,  -12'd174,  12'd154,  12'd82,  -12'd162,  -12'd171,  12'd72,  -12'd143,  
-12'd1,  12'd45,  12'd7,  12'd226,  -12'd14,  12'd261,  -12'd350,  12'd85,  -12'd342,  12'd18,  -12'd29,  12'd249,  -12'd88,  -12'd32,  -12'd191,  12'd398,  
-12'd283,  12'd130,  -12'd158,  12'd502,  12'd265,  12'd297,  12'd356,  -12'd198,  -12'd198,  -12'd0,  12'd146,  -12'd119,  -12'd9,  12'd567,  12'd136,  12'd175,  
-12'd411,  -12'd612,  -12'd78,  -12'd353,  12'd127,  -12'd225,  12'd173,  12'd197,  -12'd237,  12'd102,  -12'd121,  -12'd366,  -12'd341,  12'd231,  -12'd218,  12'd54,  
12'd105,  12'd276,  12'd182,  12'd39,  -12'd101,  -12'd101,  -12'd3,  12'd265,  -12'd116,  -12'd355,  12'd365,  12'd96,  -12'd388,  12'd260,  -12'd305,  -12'd240,  
12'd91,  -12'd4,  -12'd413,  -12'd356,  12'd76,  -12'd280,  12'd359,  -12'd113,  -12'd169,  12'd219,  -12'd16,  12'd321,  12'd47,  12'd121,  12'd302,  12'd319,  
12'd153,  12'd192,  12'd206,  12'd350,  -12'd105,  12'd134,  12'd71,  12'd177,  -12'd41,  12'd181,  12'd129,  12'd308,  12'd286,  12'd76,  12'd43,  -12'd18,  
12'd52,  -12'd131,  12'd230,  12'd78,  12'd16,  12'd249,  12'd245,  -12'd193,  -12'd10,  -12'd630,  12'd37,  12'd181,  -12'd256,  -12'd91,  12'd318,  -12'd20,  
-12'd369,  -12'd348,  12'd470,  12'd211,  12'd80,  12'd130,  12'd14,  -12'd200,  -12'd373,  -12'd35,  -12'd74,  12'd246,  -12'd142,  -12'd63,  -12'd236,  -12'd201,  
-12'd100,  12'd140,  12'd268,  -12'd409,  -12'd359,  12'd96,  12'd343,  -12'd124,  -12'd183,  -12'd30,  12'd168,  12'd66,  -12'd157,  12'd142,  -12'd89,  12'd214,  
-12'd12,  12'd107,  -12'd97,  -12'd237,  12'd3,  -12'd123,  12'd382,  -12'd124,  12'd145,  -12'd189,  12'd94,  12'd30,  12'd185,  -12'd125,  12'd111,  12'd31,  
12'd88,  12'd28,  12'd243,  12'd184,  -12'd244,  -12'd44,  12'd81,  12'd369,  12'd18,  -12'd180,  12'd87,  -12'd90,  12'd5,  12'd63,  -12'd103,  12'd27,  
12'd151,  12'd116,  12'd274,  -12'd25,  -12'd240,  -12'd69,  12'd328,  12'd317,  12'd297,  -12'd590,  12'd460,  -12'd90,  12'd312,  -12'd452,  -12'd191,  -12'd65,  
12'd294,  12'd119,  -12'd124,  -12'd187,  -12'd148,  -12'd14,  -12'd102,  12'd304,  -12'd454,  -12'd705,  -12'd18,  12'd32,  12'd213,  12'd296,  12'd451,  12'd222,  
-12'd70,  -12'd395,  -12'd320,  -12'd346,  -12'd217,  -12'd435,  12'd432,  12'd57,  -12'd264,  12'd231,  12'd69,  -12'd205,  -12'd139,  12'd33,  12'd51,  -12'd29,  
-12'd132,  12'd78,  12'd254,  -12'd59,  -12'd39,  12'd260,  12'd620,  12'd263,  12'd133,  12'd283,  -12'd112,  12'd97,  12'd142,  12'd262,  -12'd177,  -12'd121,  
-12'd173,  12'd267,  12'd475,  -12'd497,  12'd337,  -12'd638,  12'd123,  12'd191,  12'd305,  -12'd55,  -12'd206,  -12'd433,  -12'd249,  12'd131,  12'd341,  -12'd255,  
12'd45,  -12'd191,  -12'd196,  -12'd95,  -12'd221,  -12'd475,  -12'd11,  12'd103,  -12'd150,  -12'd420,  -12'd360,  -12'd537,  -12'd507,  -12'd39,  -12'd344,  -12'd93,  
-12'd173,  -12'd146,  12'd246,  -12'd254,  -12'd487,  -12'd198,  -12'd8,  12'd134,  -12'd197,  -12'd282,  -12'd270,  -12'd334,  -12'd314,  -12'd312,  -12'd205,  -12'd388,  

-12'd127,  -12'd233,  12'd95,  12'd50,  12'd33,  -12'd38,  -12'd411,  12'd418,  12'd33,  12'd267,  -12'd110,  -12'd181,  -12'd80,  -12'd59,  12'd451,  12'd392,  
-12'd130,  -12'd327,  12'd93,  12'd217,  12'd44,  12'd101,  -12'd401,  12'd140,  -12'd224,  12'd357,  12'd391,  12'd54,  12'd336,  -12'd240,  12'd219,  12'd80,  
12'd212,  -12'd5,  -12'd85,  12'd134,  12'd49,  12'd63,  12'd30,  -12'd165,  -12'd406,  12'd26,  12'd204,  12'd39,  12'd166,  -12'd920,  -12'd348,  12'd277,  
12'd387,  -12'd11,  -12'd78,  12'd54,  -12'd78,  12'd356,  12'd208,  -12'd62,  12'd331,  -12'd183,  12'd168,  12'd217,  -12'd101,  -12'd355,  -12'd104,  -12'd42,  
12'd271,  -12'd354,  12'd374,  -12'd73,  -12'd0,  -12'd101,  12'd161,  -12'd147,  12'd95,  12'd139,  -12'd147,  -12'd14,  -12'd293,  -12'd81,  -12'd235,  12'd111,  
-12'd128,  12'd162,  -12'd71,  -12'd49,  12'd286,  12'd216,  -12'd262,  12'd185,  12'd295,  -12'd92,  12'd114,  12'd183,  12'd352,  12'd5,  12'd15,  -12'd270,  
-12'd265,  -12'd225,  -12'd442,  12'd357,  12'd102,  -12'd194,  -12'd412,  -12'd137,  -12'd307,  -12'd92,  12'd145,  12'd208,  12'd331,  -12'd133,  12'd115,  -12'd144,  
12'd262,  -12'd168,  -12'd347,  12'd317,  12'd259,  12'd100,  -12'd359,  12'd286,  -12'd159,  12'd77,  12'd53,  12'd34,  12'd108,  -12'd107,  12'd87,  12'd260,  
12'd186,  12'd84,  -12'd351,  12'd100,  12'd161,  12'd52,  12'd367,  12'd367,  12'd221,  12'd198,  12'd445,  -12'd183,  12'd157,  12'd22,  -12'd36,  12'd138,  
12'd45,  -12'd559,  -12'd160,  12'd91,  -12'd262,  12'd105,  -12'd270,  12'd282,  12'd200,  12'd275,  12'd80,  -12'd95,  12'd269,  -12'd32,  -12'd90,  -12'd126,  
-12'd263,  12'd320,  -12'd112,  12'd244,  12'd276,  -12'd175,  12'd53,  12'd114,  12'd625,  12'd134,  12'd316,  12'd100,  -12'd13,  12'd232,  -12'd1,  12'd21,  
-12'd218,  -12'd50,  -12'd117,  12'd147,  12'd12,  -12'd451,  -12'd437,  -12'd196,  -12'd355,  -12'd60,  12'd277,  -12'd24,  12'd330,  -12'd112,  -12'd21,  12'd201,  
-12'd3,  -12'd161,  12'd311,  12'd77,  -12'd396,  12'd353,  12'd231,  12'd55,  -12'd232,  12'd473,  12'd157,  12'd214,  12'd153,  -12'd363,  -12'd175,  12'd331,  
12'd109,  12'd171,  -12'd338,  12'd0,  12'd182,  12'd387,  -12'd87,  12'd302,  -12'd91,  -12'd162,  -12'd74,  12'd150,  12'd37,  12'd48,  12'd138,  12'd76,  
-12'd332,  -12'd140,  -12'd207,  -12'd8,  12'd351,  -12'd169,  -12'd160,  -12'd27,  12'd75,  -12'd49,  12'd271,  12'd113,  12'd365,  12'd13,  12'd198,  -12'd306,  
-12'd74,  12'd76,  -12'd288,  -12'd345,  12'd131,  -12'd50,  -12'd182,  12'd65,  12'd277,  -12'd9,  12'd160,  12'd96,  -12'd95,  -12'd271,  -12'd447,  -12'd200,  
-12'd500,  -12'd345,  12'd175,  12'd145,  -12'd204,  -12'd235,  -12'd120,  -12'd369,  12'd36,  12'd169,  -12'd3,  12'd39,  -12'd247,  -12'd358,  12'd52,  12'd390,  
-12'd373,  12'd65,  -12'd16,  12'd61,  12'd80,  -12'd105,  12'd37,  -12'd202,  12'd443,  -12'd1,  12'd56,  12'd61,  12'd132,  -12'd457,  -12'd112,  -12'd145,  
-12'd68,  12'd180,  12'd171,  -12'd353,  -12'd284,  12'd222,  -12'd25,  -12'd120,  -12'd115,  12'd190,  12'd11,  12'd76,  -12'd1,  -12'd298,  -12'd323,  -12'd97,  
12'd223,  -12'd144,  -12'd167,  12'd96,  -12'd54,  -12'd101,  -12'd221,  12'd501,  -12'd211,  12'd158,  -12'd65,  12'd42,  12'd222,  12'd164,  -12'd73,  12'd129,  
12'd184,  12'd282,  -12'd188,  -12'd106,  12'd370,  12'd214,  12'd312,  -12'd446,  12'd238,  12'd251,  -12'd56,  12'd31,  12'd82,  -12'd226,  -12'd300,  12'd74,  
-12'd100,  -12'd166,  12'd82,  -12'd357,  -12'd103,  12'd262,  12'd292,  -12'd62,  12'd212,  12'd417,  -12'd191,  -12'd221,  -12'd112,  12'd248,  -12'd118,  12'd201,  
12'd31,  12'd411,  12'd216,  -12'd41,  -12'd139,  12'd14,  12'd459,  -12'd93,  12'd122,  12'd282,  -12'd109,  -12'd212,  12'd109,  -12'd177,  12'd190,  12'd5,  
12'd23,  -12'd310,  12'd31,  -12'd173,  12'd102,  12'd39,  12'd22,  -12'd68,  12'd200,  -12'd173,  -12'd318,  -12'd532,  -12'd557,  12'd285,  12'd36,  12'd118,  
12'd122,  -12'd134,  12'd267,  -12'd298,  -12'd105,  -12'd163,  -12'd192,  -12'd221,  12'd158,  -12'd209,  -12'd75,  -12'd108,  12'd102,  -12'd312,  -12'd280,  12'd19,  

12'd397,  12'd42,  12'd35,  -12'd14,  -12'd115,  -12'd241,  12'd192,  12'd8,  12'd105,  -12'd116,  -12'd137,  -12'd147,  12'd5,  12'd37,  -12'd473,  -12'd204,  
12'd560,  12'd77,  12'd271,  -12'd64,  -12'd9,  12'd153,  12'd323,  -12'd16,  12'd51,  -12'd26,  12'd215,  12'd132,  12'd20,  12'd100,  -12'd123,  12'd401,  
12'd478,  12'd27,  12'd37,  12'd308,  -12'd80,  -12'd296,  12'd92,  12'd139,  -12'd99,  -12'd62,  12'd205,  12'd22,  12'd379,  -12'd227,  12'd76,  12'd91,  
-12'd217,  12'd210,  12'd395,  12'd79,  -12'd34,  12'd248,  -12'd612,  -12'd217,  -12'd408,  -12'd102,  -12'd144,  -12'd253,  12'd188,  -12'd140,  12'd44,  -12'd136,  
12'd113,  -12'd103,  12'd50,  -12'd12,  12'd418,  -12'd312,  -12'd109,  -12'd275,  -12'd534,  -12'd191,  -12'd62,  -12'd279,  12'd330,  12'd96,  12'd5,  12'd633,  
12'd323,  -12'd422,  12'd379,  -12'd63,  -12'd13,  12'd352,  -12'd78,  12'd249,  -12'd10,  -12'd42,  -12'd311,  -12'd213,  12'd17,  12'd137,  12'd51,  -12'd258,  
-12'd53,  -12'd253,  -12'd33,  -12'd136,  -12'd69,  -12'd25,  -12'd83,  -12'd117,  -12'd218,  12'd10,  12'd95,  12'd309,  -12'd250,  -12'd168,  -12'd7,  -12'd158,  
-12'd73,  12'd113,  -12'd208,  -12'd226,  12'd320,  12'd191,  12'd16,  12'd87,  12'd251,  12'd450,  12'd287,  -12'd33,  -12'd88,  -12'd154,  -12'd68,  12'd80,  
-12'd95,  -12'd20,  -12'd72,  -12'd94,  12'd121,  -12'd272,  -12'd464,  12'd94,  -12'd210,  12'd517,  12'd267,  -12'd80,  12'd55,  -12'd331,  -12'd271,  12'd198,  
-12'd144,  -12'd49,  -12'd154,  -12'd141,  12'd465,  12'd237,  -12'd222,  12'd169,  -12'd93,  12'd145,  12'd93,  12'd45,  -12'd22,  12'd47,  -12'd188,  12'd192,  
12'd52,  12'd9,  12'd44,  -12'd132,  12'd214,  -12'd3,  -12'd226,  -12'd109,  -12'd279,  12'd144,  -12'd319,  12'd107,  -12'd314,  12'd91,  12'd353,  -12'd107,  
-12'd168,  12'd65,  -12'd137,  12'd57,  12'd254,  12'd241,  -12'd170,  -12'd228,  12'd55,  12'd71,  12'd16,  12'd15,  -12'd180,  -12'd279,  12'd37,  -12'd46,  
12'd75,  -12'd207,  12'd75,  12'd331,  12'd229,  12'd26,  -12'd24,  12'd319,  12'd478,  -12'd47,  -12'd51,  12'd110,  -12'd484,  -12'd113,  -12'd88,  12'd11,  
12'd356,  -12'd159,  -12'd158,  -12'd93,  -12'd137,  12'd98,  -12'd165,  -12'd46,  12'd225,  12'd644,  12'd44,  -12'd151,  12'd234,  12'd109,  -12'd528,  12'd66,  
12'd152,  12'd149,  -12'd302,  -12'd110,  12'd397,  12'd167,  -12'd84,  -12'd241,  12'd121,  12'd403,  12'd163,  12'd234,  -12'd199,  -12'd1,  -12'd213,  -12'd60,  
12'd248,  12'd117,  -12'd104,  12'd268,  -12'd31,  -12'd341,  12'd106,  -12'd63,  -12'd243,  12'd219,  -12'd365,  12'd149,  12'd18,  12'd187,  12'd101,  12'd127,  
12'd399,  12'd369,  12'd139,  12'd415,  -12'd11,  -12'd79,  12'd18,  -12'd152,  12'd350,  12'd357,  -12'd31,  12'd271,  -12'd119,  12'd170,  12'd116,  -12'd308,  
12'd259,  12'd319,  -12'd17,  12'd99,  12'd349,  12'd59,  -12'd295,  -12'd89,  -12'd173,  -12'd116,  12'd243,  12'd86,  -12'd137,  12'd213,  -12'd54,  12'd208,  
-12'd194,  12'd212,  -12'd256,  -12'd86,  12'd155,  -12'd375,  -12'd246,  12'd54,  -12'd237,  -12'd93,  -12'd55,  -12'd40,  12'd57,  -12'd86,  12'd502,  -12'd178,  
12'd4,  -12'd112,  12'd182,  -12'd44,  -12'd417,  12'd340,  -12'd344,  12'd296,  12'd122,  12'd21,  -12'd12,  12'd262,  12'd279,  12'd206,  -12'd28,  12'd72,  
12'd308,  12'd17,  12'd75,  12'd183,  -12'd309,  12'd192,  12'd0,  12'd308,  12'd232,  12'd307,  -12'd7,  12'd173,  12'd7,  12'd593,  -12'd11,  -12'd118,  
12'd82,  12'd56,  12'd35,  12'd293,  12'd226,  12'd22,  -12'd195,  12'd240,  12'd56,  -12'd103,  12'd202,  -12'd152,  12'd169,  12'd214,  12'd504,  -12'd49,  
-12'd166,  -12'd108,  -12'd343,  12'd12,  12'd250,  12'd149,  -12'd170,  12'd62,  -12'd142,  -12'd343,  -12'd55,  -12'd48,  12'd230,  -12'd663,  12'd130,  -12'd26,  
12'd152,  12'd58,  12'd88,  -12'd57,  12'd81,  12'd324,  12'd17,  12'd440,  12'd49,  -12'd82,  -12'd105,  12'd322,  12'd167,  12'd49,  -12'd19,  12'd140,  
12'd83,  12'd217,  12'd312,  -12'd0,  -12'd201,  12'd77,  12'd239,  12'd169,  12'd345,  12'd113,  -12'd282,  12'd551,  -12'd214,  -12'd111,  12'd2,  12'd2,  

-12'd247,  12'd202,  -12'd161,  12'd115,  12'd446,  -12'd59,  -12'd356,  12'd198,  -12'd253,  12'd81,  -12'd50,  12'd57,  -12'd41,  12'd221,  -12'd57,  12'd515,  
-12'd281,  12'd201,  12'd83,  12'd252,  12'd165,  12'd222,  -12'd173,  -12'd46,  12'd123,  12'd249,  -12'd348,  12'd192,  -12'd84,  -12'd391,  12'd463,  12'd598,  
-12'd238,  -12'd35,  12'd279,  12'd129,  -12'd72,  -12'd229,  12'd46,  12'd143,  12'd15,  12'd18,  -12'd252,  12'd88,  12'd182,  12'd217,  -12'd305,  12'd303,  
-12'd126,  -12'd423,  12'd31,  -12'd4,  12'd44,  -12'd124,  12'd353,  -12'd201,  -12'd5,  -12'd162,  12'd141,  12'd296,  -12'd288,  12'd681,  12'd34,  -12'd426,  
-12'd372,  12'd155,  12'd274,  -12'd282,  -12'd287,  -12'd122,  12'd84,  -12'd309,  12'd69,  -12'd82,  -12'd375,  -12'd281,  -12'd405,  12'd304,  -12'd375,  -12'd276,  
12'd248,  12'd309,  -12'd208,  -12'd166,  12'd172,  -12'd82,  -12'd126,  12'd169,  -12'd82,  -12'd285,  12'd87,  12'd12,  12'd98,  -12'd279,  12'd203,  12'd278,  
12'd36,  12'd120,  -12'd196,  -12'd227,  12'd72,  12'd167,  -12'd106,  -12'd153,  12'd41,  12'd511,  12'd199,  12'd293,  -12'd82,  12'd7,  12'd268,  12'd94,  
12'd474,  12'd141,  12'd483,  12'd176,  -12'd268,  -12'd188,  12'd22,  -12'd12,  12'd47,  12'd139,  -12'd68,  12'd322,  12'd38,  -12'd224,  12'd43,  12'd5,  
12'd387,  -12'd198,  12'd159,  12'd339,  12'd15,  12'd379,  12'd445,  -12'd59,  -12'd263,  12'd198,  12'd83,  12'd137,  12'd39,  12'd736,  -12'd136,  -12'd132,  
12'd228,  -12'd77,  12'd67,  12'd105,  12'd306,  12'd364,  12'd53,  -12'd415,  -12'd0,  -12'd281,  12'd100,  -12'd133,  12'd119,  12'd441,  -12'd453,  -12'd331,  
-12'd547,  -12'd112,  -12'd258,  12'd8,  12'd6,  -12'd242,  12'd199,  12'd99,  12'd341,  12'd130,  -12'd68,  -12'd198,  -12'd122,  -12'd163,  -12'd443,  12'd142,  
12'd167,  12'd31,  -12'd7,  12'd12,  -12'd91,  -12'd69,  -12'd331,  12'd317,  -12'd241,  12'd1,  -12'd89,  -12'd176,  12'd187,  12'd374,  12'd157,  12'd5,  
12'd176,  -12'd211,  -12'd243,  -12'd48,  12'd28,  -12'd88,  -12'd50,  12'd287,  -12'd687,  12'd106,  12'd224,  -12'd88,  12'd351,  -12'd86,  12'd192,  -12'd245,  
-12'd0,  -12'd150,  12'd224,  12'd384,  12'd100,  12'd169,  -12'd66,  12'd197,  -12'd116,  12'd117,  12'd318,  12'd115,  12'd197,  -12'd141,  -12'd235,  12'd47,  
-12'd149,  -12'd394,  -12'd27,  -12'd354,  12'd249,  12'd62,  -12'd31,  12'd125,  -12'd34,  12'd93,  12'd133,  12'd100,  12'd368,  12'd31,  -12'd273,  -12'd50,  
-12'd594,  -12'd499,  12'd91,  12'd210,  12'd208,  -12'd0,  -12'd379,  12'd294,  12'd296,  -12'd28,  12'd12,  -12'd518,  -12'd177,  -12'd51,  -12'd111,  -12'd245,  
-12'd296,  12'd45,  12'd165,  -12'd127,  12'd104,  12'd69,  -12'd185,  -12'd271,  -12'd73,  12'd159,  12'd97,  -12'd239,  -12'd148,  -12'd354,  -12'd22,  -12'd72,  
-12'd239,  12'd224,  12'd72,  -12'd162,  -12'd263,  -12'd155,  -12'd74,  12'd198,  12'd79,  12'd214,  12'd239,  12'd41,  -12'd336,  -12'd130,  12'd46,  12'd55,  
-12'd194,  -12'd59,  -12'd18,  -12'd334,  -12'd159,  12'd226,  -12'd181,  12'd83,  12'd107,  -12'd218,  12'd243,  -12'd151,  -12'd22,  12'd320,  -12'd183,  12'd46,  
12'd49,  12'd273,  12'd23,  -12'd274,  12'd102,  12'd24,  12'd50,  -12'd166,  -12'd67,  -12'd153,  12'd2,  -12'd205,  12'd237,  12'd23,  12'd57,  12'd111,  
-12'd304,  -12'd312,  -12'd81,  -12'd18,  12'd76,  -12'd84,  12'd507,  -12'd223,  -12'd21,  -12'd11,  -12'd161,  12'd269,  12'd382,  -12'd202,  12'd212,  -12'd106,  
12'd472,  -12'd71,  12'd132,  -12'd137,  12'd309,  12'd57,  12'd251,  -12'd282,  12'd159,  -12'd53,  -12'd18,  12'd253,  -12'd179,  -12'd8,  12'd197,  12'd202,  
12'd198,  12'd401,  12'd145,  12'd12,  12'd58,  12'd99,  12'd47,  12'd58,  -12'd108,  -12'd210,  -12'd21,  12'd215,  12'd25,  12'd146,  -12'd237,  12'd78,  
-12'd122,  -12'd131,  12'd99,  -12'd195,  -12'd135,  -12'd332,  12'd294,  12'd27,  -12'd228,  12'd100,  12'd161,  12'd92,  -12'd36,  12'd242,  -12'd108,  12'd36,  
12'd192,  12'd214,  12'd223,  12'd211,  12'd184,  -12'd450,  12'd381,  -12'd147,  -12'd60,  12'd127,  12'd37,  12'd160,  -12'd164,  12'd187,  -12'd154,  -12'd187,  

-12'd52,  -12'd59,  -12'd128,  -12'd93,  -12'd304,  12'd94,  -12'd437,  -12'd18,  -12'd479,  -12'd165,  12'd490,  -12'd190,  -12'd2,  -12'd340,  12'd123,  12'd128,  
-12'd6,  12'd140,  -12'd434,  12'd181,  12'd364,  12'd299,  -12'd197,  12'd305,  12'd339,  -12'd53,  -12'd55,  12'd306,  12'd148,  -12'd355,  12'd147,  -12'd91,  
-12'd62,  12'd240,  12'd205,  -12'd71,  12'd166,  12'd205,  -12'd416,  12'd157,  12'd214,  -12'd305,  -12'd188,  12'd245,  12'd148,  -12'd453,  12'd133,  12'd151,  
12'd198,  -12'd78,  12'd396,  12'd37,  -12'd121,  12'd69,  12'd280,  12'd289,  12'd113,  12'd397,  12'd165,  -12'd60,  12'd486,  -12'd242,  12'd118,  12'd47,  
-12'd122,  -12'd694,  -12'd114,  12'd39,  -12'd105,  12'd277,  12'd191,  -12'd114,  -12'd100,  12'd313,  12'd242,  -12'd254,  -12'd147,  -12'd224,  12'd21,  -12'd109,  
-12'd170,  -12'd301,  12'd5,  -12'd248,  12'd21,  -12'd84,  12'd63,  -12'd337,  -12'd174,  -12'd384,  12'd139,  -12'd216,  -12'd170,  12'd14,  -12'd207,  12'd89,  
12'd6,  12'd36,  -12'd426,  12'd49,  -12'd23,  12'd235,  12'd137,  -12'd227,  -12'd108,  12'd210,  -12'd60,  -12'd134,  12'd27,  -12'd42,  -12'd461,  12'd303,  
-12'd292,  12'd464,  -12'd173,  -12'd284,  -12'd60,  12'd39,  12'd65,  -12'd119,  12'd44,  12'd172,  12'd97,  -12'd204,  12'd65,  12'd485,  -12'd233,  -12'd110,  
12'd114,  12'd185,  12'd54,  -12'd61,  12'd11,  12'd417,  12'd365,  -12'd104,  12'd249,  -12'd167,  -12'd179,  12'd285,  -12'd17,  12'd617,  12'd264,  12'd23,  
-12'd605,  12'd459,  12'd338,  12'd94,  12'd111,  -12'd70,  -12'd200,  -12'd247,  -12'd40,  -12'd413,  12'd108,  -12'd417,  -12'd542,  12'd188,  12'd556,  -12'd233,  
-12'd313,  -12'd243,  -12'd252,  -12'd55,  -12'd245,  -12'd441,  12'd280,  -12'd259,  -12'd188,  12'd158,  12'd75,  12'd72,  -12'd268,  -12'd252,  12'd48,  -12'd194,  
-12'd26,  12'd25,  -12'd243,  12'd14,  -12'd20,  12'd61,  12'd156,  -12'd249,  12'd378,  -12'd27,  -12'd277,  12'd220,  12'd121,  -12'd760,  -12'd76,  12'd93,  
-12'd81,  12'd55,  -12'd163,  -12'd361,  -12'd3,  -12'd322,  12'd230,  -12'd94,  12'd80,  12'd238,  -12'd25,  -12'd187,  -12'd58,  12'd173,  -12'd35,  -12'd15,  
12'd185,  12'd82,  12'd170,  12'd332,  -12'd160,  12'd86,  12'd85,  -12'd64,  12'd17,  -12'd484,  -12'd170,  12'd391,  -12'd141,  12'd57,  12'd136,  -12'd488,  
12'd470,  -12'd40,  -12'd92,  12'd336,  -12'd448,  12'd120,  -12'd88,  -12'd6,  -12'd49,  -12'd84,  -12'd22,  12'd264,  -12'd40,  12'd72,  12'd226,  -12'd400,  
12'd281,  -12'd272,  12'd240,  12'd228,  -12'd690,  12'd20,  12'd368,  -12'd3,  12'd177,  12'd80,  12'd262,  12'd9,  -12'd135,  -12'd41,  -12'd25,  12'd149,  
12'd20,  -12'd428,  -12'd32,  -12'd90,  -12'd344,  -12'd76,  -12'd224,  -12'd4,  12'd121,  12'd155,  -12'd140,  12'd389,  12'd348,  -12'd143,  -12'd139,  12'd4,  
12'd277,  -12'd228,  12'd153,  -12'd54,  -12'd175,  12'd286,  -12'd154,  12'd217,  -12'd68,  -12'd123,  -12'd474,  12'd113,  12'd251,  12'd151,  12'd207,  -12'd52,  
12'd143,  12'd27,  12'd120,  12'd261,  -12'd40,  12'd171,  12'd187,  12'd298,  12'd422,  12'd348,  -12'd147,  12'd27,  -12'd23,  -12'd274,  -12'd177,  -12'd136,  
12'd276,  12'd184,  -12'd441,  12'd143,  -12'd15,  12'd181,  12'd38,  12'd189,  -12'd9,  12'd227,  12'd329,  12'd37,  12'd132,  12'd128,  12'd115,  12'd92,  
12'd82,  -12'd180,  12'd332,  -12'd235,  -12'd181,  12'd138,  -12'd5,  12'd38,  -12'd186,  -12'd36,  12'd79,  -12'd80,  -12'd45,  12'd206,  -12'd81,  12'd266,  
-12'd138,  12'd164,  -12'd350,  -12'd101,  -12'd40,  12'd265,  12'd212,  -12'd4,  12'd230,  -12'd340,  12'd257,  -12'd250,  12'd104,  12'd90,  12'd202,  12'd72,  
-12'd125,  12'd278,  12'd137,  -12'd94,  -12'd146,  -12'd181,  -12'd195,  12'd133,  -12'd247,  -12'd226,  12'd71,  -12'd219,  12'd179,  12'd305,  -12'd158,  -12'd201,  
-12'd408,  12'd150,  -12'd6,  12'd177,  -12'd40,  12'd115,  -12'd83,  12'd117,  -12'd209,  -12'd51,  -12'd11,  -12'd275,  12'd24,  12'd94,  12'd60,  12'd58,  
-12'd68,  -12'd172,  -12'd509,  -12'd176,  -12'd107,  12'd121,  12'd150,  12'd74,  -12'd580,  12'd839,  12'd160,  12'd75,  -12'd160,  -12'd112,  -12'd176,  12'd283,  

-12'd184,  -12'd126,  12'd157,  -12'd234,  -12'd34,  -12'd182,  12'd822,  -12'd232,  12'd302,  12'd100,  12'd149,  12'd37,  -12'd35,  12'd141,  12'd300,  12'd405,  
-12'd345,  12'd118,  12'd199,  -12'd354,  -12'd472,  12'd130,  12'd728,  12'd30,  -12'd336,  12'd22,  12'd177,  12'd195,  12'd277,  12'd432,  -12'd157,  -12'd50,  
12'd163,  -12'd113,  12'd258,  -12'd458,  -12'd55,  -12'd175,  12'd455,  -12'd10,  -12'd362,  -12'd451,  12'd156,  12'd274,  -12'd434,  12'd477,  -12'd141,  -12'd714,  
12'd744,  12'd133,  -12'd395,  -12'd252,  -12'd85,  12'd21,  12'd363,  -12'd129,  -12'd259,  -12'd296,  -12'd12,  12'd86,  12'd44,  12'd257,  -12'd391,  -12'd310,  
12'd205,  12'd350,  -12'd116,  -12'd25,  -12'd438,  -12'd120,  12'd28,  -12'd177,  12'd100,  12'd14,  -12'd131,  -12'd174,  -12'd370,  -12'd12,  12'd51,  12'd73,  
12'd255,  -12'd167,  12'd254,  -12'd15,  12'd41,  -12'd344,  12'd633,  -12'd291,  -12'd96,  12'd191,  12'd437,  -12'd184,  12'd40,  -12'd184,  12'd113,  12'd283,  
-12'd256,  12'd145,  12'd24,  -12'd61,  12'd261,  -12'd150,  12'd342,  -12'd368,  -12'd223,  -12'd178,  12'd310,  12'd38,  12'd92,  -12'd116,  -12'd549,  -12'd90,  
12'd489,  12'd288,  12'd224,  -12'd264,  -12'd417,  12'd0,  -12'd267,  -12'd99,  -12'd81,  12'd122,  -12'd201,  12'd14,  12'd261,  12'd117,  12'd86,  12'd34,  
12'd404,  12'd461,  -12'd145,  12'd166,  -12'd88,  12'd346,  -12'd209,  -12'd212,  12'd275,  12'd214,  12'd71,  12'd138,  12'd87,  12'd134,  12'd34,  12'd23,  
-12'd4,  -12'd323,  12'd103,  12'd232,  12'd189,  -12'd418,  -12'd77,  -12'd33,  -12'd1,  -12'd7,  12'd36,  12'd326,  12'd261,  -12'd330,  12'd231,  12'd86,  
12'd54,  -12'd366,  -12'd7,  -12'd65,  -12'd107,  -12'd243,  12'd702,  -12'd108,  -12'd127,  -12'd198,  12'd74,  12'd317,  -12'd519,  -12'd552,  12'd234,  -12'd330,  
12'd363,  -12'd355,  -12'd259,  -12'd156,  -12'd139,  12'd278,  -12'd282,  -12'd105,  12'd241,  -12'd346,  12'd99,  12'd50,  -12'd261,  -12'd40,  -12'd45,  12'd41,  
12'd380,  12'd141,  -12'd13,  -12'd108,  -12'd60,  -12'd232,  -12'd3,  -12'd50,  -12'd61,  -12'd55,  -12'd488,  -12'd147,  12'd178,  -12'd296,  -12'd94,  -12'd144,  
-12'd8,  12'd250,  -12'd200,  -12'd206,  -12'd44,  12'd336,  12'd81,  -12'd245,  12'd161,  12'd307,  -12'd82,  12'd128,  -12'd27,  12'd19,  -12'd50,  -12'd90,  
-12'd144,  -12'd45,  12'd176,  12'd357,  -12'd159,  12'd71,  -12'd23,  -12'd31,  -12'd181,  12'd120,  -12'd382,  12'd198,  12'd186,  -12'd14,  12'd222,  12'd0,  
12'd119,  12'd73,  12'd136,  12'd56,  12'd185,  12'd133,  12'd338,  12'd243,  -12'd29,  12'd69,  -12'd218,  12'd147,  -12'd47,  12'd59,  -12'd36,  12'd5,  
12'd6,  -12'd181,  12'd81,  12'd329,  12'd40,  -12'd170,  12'd60,  -12'd344,  12'd88,  12'd34,  12'd168,  -12'd151,  12'd103,  12'd210,  -12'd10,  12'd134,  
12'd169,  -12'd250,  12'd20,  12'd142,  -12'd441,  -12'd142,  -12'd260,  12'd347,  12'd232,  12'd345,  -12'd184,  -12'd172,  12'd391,  -12'd245,  12'd53,  -12'd1,  
12'd389,  -12'd288,  -12'd297,  12'd84,  -12'd370,  -12'd109,  -12'd249,  12'd183,  -12'd162,  -12'd96,  12'd358,  12'd47,  12'd471,  12'd225,  12'd111,  -12'd352,  
12'd59,  -12'd43,  12'd211,  12'd144,  -12'd13,  -12'd176,  12'd153,  12'd197,  12'd92,  12'd267,  -12'd197,  -12'd17,  12'd499,  -12'd99,  -12'd48,  12'd194,  
-12'd149,  12'd168,  12'd3,  12'd446,  12'd156,  12'd346,  -12'd242,  12'd95,  12'd315,  12'd125,  12'd175,  -12'd414,  -12'd72,  -12'd206,  -12'd68,  12'd123,  
12'd39,  -12'd205,  12'd7,  12'd97,  -12'd100,  -12'd343,  12'd275,  -12'd155,  12'd122,  12'd228,  12'd36,  -12'd325,  12'd236,  -12'd220,  -12'd187,  12'd49,  
-12'd147,  12'd32,  -12'd216,  12'd6,  -12'd240,  12'd126,  -12'd17,  -12'd134,  -12'd40,  12'd444,  -12'd90,  12'd30,  12'd245,  -12'd338,  12'd102,  12'd352,  
-12'd584,  -12'd195,  -12'd204,  12'd90,  12'd49,  12'd268,  -12'd175,  -12'd367,  -12'd161,  12'd278,  -12'd195,  -12'd245,  -12'd171,  -12'd168,  -12'd406,  12'd220,  
-12'd144,  -12'd24,  -12'd92,  -12'd94,  12'd110,  -12'd262,  -12'd418,  12'd67,  -12'd104,  -12'd153,  12'd238,  -12'd307,  12'd39,  -12'd30,  -12'd70,  -12'd43,  

-12'd125,  -12'd459,  -12'd33,  12'd175,  12'd200,  -12'd41,  -12'd358,  12'd90,  -12'd78,  12'd58,  12'd199,  -12'd47,  -12'd84,  -12'd166,  -12'd118,  -12'd464,  
-12'd55,  -12'd181,  -12'd412,  12'd334,  -12'd96,  12'd215,  -12'd172,  12'd392,  12'd56,  12'd306,  -12'd1,  -12'd138,  -12'd165,  -12'd236,  12'd300,  -12'd267,  
-12'd116,  -12'd29,  12'd66,  12'd380,  -12'd252,  12'd110,  -12'd183,  -12'd67,  -12'd69,  12'd100,  -12'd199,  -12'd55,  12'd251,  12'd151,  12'd321,  12'd258,  
12'd5,  -12'd132,  12'd307,  12'd35,  -12'd67,  -12'd121,  -12'd2,  12'd315,  -12'd30,  12'd360,  12'd107,  -12'd335,  -12'd178,  -12'd664,  12'd305,  12'd336,  
12'd116,  12'd115,  12'd380,  -12'd28,  12'd59,  12'd191,  -12'd348,  12'd293,  12'd132,  -12'd81,  -12'd367,  12'd192,  12'd201,  12'd151,  12'd321,  -12'd336,  
-12'd216,  -12'd184,  12'd2,  -12'd93,  12'd349,  12'd115,  -12'd287,  -12'd5,  12'd32,  12'd142,  -12'd219,  -12'd203,  12'd350,  12'd200,  -12'd412,  12'd160,  
12'd260,  12'd284,  12'd326,  -12'd19,  -12'd143,  12'd453,  -12'd95,  12'd30,  -12'd112,  12'd191,  12'd457,  -12'd284,  12'd63,  12'd101,  12'd153,  12'd48,  
-12'd422,  12'd484,  12'd87,  -12'd1,  12'd41,  12'd335,  12'd1,  -12'd145,  12'd72,  -12'd76,  -12'd172,  -12'd309,  -12'd242,  12'd226,  12'd291,  12'd170,  
-12'd552,  12'd487,  12'd314,  12'd337,  12'd364,  12'd221,  -12'd500,  12'd236,  -12'd8,  -12'd99,  12'd46,  -12'd289,  -12'd153,  -12'd191,  12'd164,  12'd83,  
12'd211,  12'd315,  12'd296,  12'd187,  -12'd183,  12'd438,  12'd274,  12'd115,  -12'd30,  -12'd103,  -12'd8,  -12'd66,  -12'd139,  12'd28,  12'd321,  12'd199,  
-12'd251,  -12'd158,  12'd90,  -12'd378,  -12'd126,  -12'd202,  -12'd376,  -12'd156,  -12'd65,  -12'd27,  -12'd203,  12'd104,  -12'd11,  -12'd127,  -12'd169,  -12'd76,  
12'd181,  -12'd192,  12'd79,  -12'd155,  12'd117,  12'd191,  12'd71,  -12'd34,  -12'd40,  -12'd120,  12'd248,  -12'd25,  -12'd250,  12'd315,  12'd229,  12'd249,  
12'd28,  12'd7,  -12'd91,  -12'd50,  12'd235,  12'd136,  12'd184,  12'd272,  -12'd117,  -12'd234,  -12'd151,  -12'd123,  -12'd73,  12'd58,  -12'd75,  -12'd114,  
-12'd38,  12'd325,  12'd87,  12'd91,  -12'd4,  -12'd107,  12'd48,  -12'd154,  12'd241,  -12'd1,  12'd127,  -12'd107,  -12'd113,  12'd235,  12'd437,  -12'd242,  
12'd672,  12'd331,  12'd186,  -12'd137,  12'd116,  -12'd361,  -12'd148,  -12'd182,  -12'd64,  -12'd160,  -12'd421,  -12'd25,  12'd171,  -12'd56,  12'd123,  -12'd40,  
12'd387,  -12'd8,  12'd116,  12'd79,  12'd280,  -12'd182,  12'd76,  -12'd357,  12'd295,  12'd104,  -12'd166,  12'd222,  -12'd420,  12'd100,  -12'd36,  12'd13,  
12'd441,  -12'd193,  12'd14,  -12'd31,  -12'd336,  12'd145,  12'd516,  -12'd148,  12'd295,  -12'd10,  12'd163,  12'd334,  12'd134,  12'd137,  -12'd177,  -12'd55,  
-12'd22,  -12'd319,  -12'd176,  -12'd12,  12'd338,  12'd218,  -12'd17,  -12'd81,  12'd58,  12'd260,  12'd277,  12'd6,  12'd169,  12'd429,  -12'd36,  -12'd3,  
-12'd216,  12'd31,  -12'd325,  12'd198,  12'd35,  -12'd413,  -12'd379,  -12'd163,  -12'd45,  12'd30,  -12'd334,  12'd135,  -12'd113,  -12'd248,  -12'd163,  -12'd397,  
12'd17,  -12'd36,  12'd357,  -12'd187,  12'd49,  -12'd208,  -12'd284,  -12'd180,  -12'd278,  -12'd174,  12'd193,  -12'd32,  -12'd1,  -12'd459,  -12'd96,  12'd75,  
-12'd22,  12'd37,  12'd106,  -12'd67,  12'd41,  12'd312,  -12'd329,  12'd312,  -12'd40,  -12'd15,  12'd62,  12'd59,  12'd112,  12'd277,  12'd34,  -12'd86,  
-12'd173,  12'd233,  12'd188,  12'd57,  -12'd85,  12'd100,  -12'd55,  -12'd40,  12'd134,  -12'd263,  12'd99,  12'd22,  -12'd54,  12'd394,  12'd332,  12'd129,  
12'd127,  -12'd299,  12'd265,  -12'd118,  12'd227,  12'd21,  -12'd275,  -12'd5,  -12'd166,  -12'd71,  12'd32,  -12'd16,  12'd65,  -12'd290,  12'd354,  12'd111,  
-12'd149,  -12'd231,  -12'd144,  -12'd29,  12'd62,  12'd111,  12'd52,  12'd117,  -12'd126,  -12'd392,  12'd384,  12'd217,  12'd276,  12'd125,  -12'd237,  -12'd27,  
12'd331,  -12'd89,  12'd192,  -12'd344,  -12'd318,  -12'd124,  12'd95,  12'd52,  12'd105,  -12'd420,  -12'd65,  12'd141,  -12'd234,  -12'd34,  -12'd410,  -12'd245,  

12'd41,  -12'd51,  12'd466,  -12'd93,  12'd39,  -12'd167,  12'd353,  -12'd230,  12'd244,  12'd118,  -12'd85,  -12'd154,  -12'd181,  12'd278,  -12'd139,  -12'd438,  
-12'd31,  -12'd223,  12'd9,  12'd137,  12'd60,  12'd172,  12'd687,  12'd24,  12'd21,  -12'd283,  12'd53,  12'd93,  12'd93,  12'd37,  -12'd194,  -12'd284,  
12'd135,  12'd375,  -12'd203,  -12'd30,  12'd84,  -12'd107,  -12'd73,  -12'd40,  12'd316,  -12'd248,  12'd202,  -12'd116,  12'd320,  -12'd62,  -12'd441,  -12'd223,  
12'd121,  12'd420,  -12'd212,  12'd247,  -12'd207,  12'd375,  -12'd123,  -12'd162,  -12'd71,  -12'd248,  12'd20,  12'd209,  12'd347,  -12'd115,  12'd126,  12'd293,  
12'd287,  12'd415,  -12'd30,  12'd185,  -12'd65,  -12'd186,  -12'd151,  12'd187,  -12'd367,  -12'd69,  -12'd84,  -12'd193,  12'd704,  12'd78,  12'd106,  12'd287,  
12'd258,  -12'd102,  12'd350,  12'd254,  -12'd157,  12'd25,  -12'd73,  12'd48,  12'd452,  12'd471,  -12'd347,  12'd32,  12'd605,  12'd221,  12'd415,  -12'd86,  
-12'd190,  12'd181,  12'd161,  -12'd86,  12'd61,  -12'd200,  -12'd308,  -12'd121,  12'd5,  12'd76,  -12'd8,  -12'd37,  -12'd252,  -12'd3,  12'd330,  12'd20,  
12'd47,  -12'd34,  -12'd127,  -12'd274,  -12'd210,  -12'd268,  -12'd154,  -12'd242,  12'd238,  12'd248,  12'd526,  -12'd193,  12'd2,  -12'd162,  -12'd39,  12'd101,  
-12'd348,  12'd28,  -12'd153,  -12'd133,  -12'd286,  12'd0,  -12'd103,  -12'd592,  -12'd139,  12'd132,  -12'd99,  12'd21,  12'd268,  -12'd323,  -12'd237,  12'd141,  
12'd212,  -12'd278,  -12'd319,  -12'd137,  12'd165,  12'd210,  -12'd334,  12'd136,  -12'd175,  12'd472,  12'd89,  12'd165,  12'd163,  -12'd122,  12'd124,  12'd33,  
-12'd148,  12'd366,  12'd276,  12'd384,  12'd143,  12'd123,  -12'd685,  -12'd214,  12'd2,  12'd118,  -12'd242,  -12'd66,  12'd37,  12'd483,  12'd308,  12'd47,  
-12'd102,  12'd197,  12'd1,  12'd158,  -12'd157,  -12'd36,  12'd68,  -12'd41,  -12'd203,  -12'd129,  12'd130,  12'd185,  -12'd117,  12'd300,  12'd50,  -12'd6,  
-12'd459,  -12'd327,  -12'd323,  -12'd6,  12'd212,  12'd233,  12'd139,  -12'd58,  12'd237,  -12'd600,  -12'd79,  12'd261,  -12'd42,  -12'd358,  -12'd48,  -12'd271,  
-12'd230,  12'd251,  -12'd383,  12'd154,  12'd402,  -12'd395,  -12'd98,  12'd14,  12'd169,  12'd220,  12'd41,  12'd63,  12'd38,  12'd120,  -12'd152,  -12'd16,  
-12'd290,  -12'd294,  -12'd192,  12'd152,  12'd212,  12'd317,  -12'd545,  -12'd20,  12'd49,  12'd577,  12'd103,  12'd232,  12'd224,  12'd50,  -12'd5,  -12'd190,  
-12'd60,  -12'd63,  12'd313,  -12'd74,  12'd165,  12'd31,  12'd169,  12'd149,  -12'd113,  -12'd140,  -12'd208,  12'd103,  -12'd112,  12'd147,  -12'd103,  -12'd154,  
12'd291,  12'd27,  12'd284,  -12'd36,  -12'd87,  -12'd179,  -12'd229,  12'd310,  12'd119,  12'd261,  -12'd97,  12'd402,  -12'd81,  12'd359,  12'd291,  12'd62,  
-12'd149,  12'd77,  -12'd250,  -12'd81,  12'd313,  12'd289,  12'd3,  12'd153,  -12'd207,  -12'd154,  12'd28,  12'd258,  -12'd273,  -12'd666,  12'd198,  12'd266,  
-12'd275,  -12'd93,  -12'd253,  -12'd358,  12'd359,  -12'd18,  -12'd216,  -12'd432,  12'd83,  -12'd81,  12'd223,  -12'd292,  12'd79,  12'd159,  12'd331,  12'd289,  
-12'd178,  -12'd229,  12'd577,  -12'd97,  -12'd125,  -12'd56,  -12'd47,  -12'd281,  12'd158,  -12'd237,  -12'd2,  12'd90,  -12'd10,  12'd15,  -12'd413,  -12'd192,  
12'd252,  -12'd303,  -12'd0,  -12'd270,  12'd41,  12'd134,  -12'd25,  12'd217,  12'd433,  -12'd224,  -12'd232,  12'd8,  12'd19,  12'd392,  -12'd3,  12'd8,  
12'd330,  12'd127,  12'd62,  12'd182,  12'd174,  -12'd319,  -12'd329,  -12'd87,  -12'd52,  -12'd76,  -12'd89,  -12'd1,  12'd234,  -12'd3,  12'd350,  12'd127,  
-12'd19,  -12'd39,  -12'd273,  -12'd73,  -12'd113,  12'd155,  12'd126,  12'd93,  -12'd155,  -12'd570,  -12'd11,  12'd6,  12'd149,  -12'd437,  12'd189,  12'd18,  
-12'd203,  -12'd247,  -12'd325,  -12'd360,  -12'd179,  12'd62,  -12'd130,  12'd263,  12'd261,  -12'd474,  12'd218,  12'd179,  12'd209,  12'd300,  -12'd129,  -12'd81,  
-12'd30,  12'd129,  -12'd534,  -12'd61,  -12'd260,  12'd55,  12'd113,  12'd247,  -12'd94,  -12'd926,  12'd28,  -12'd15,  -12'd136,  -12'd210,  -12'd60,  -12'd165,  

-12'd138,  12'd82,  12'd273,  -12'd78,  -12'd75,  12'd112,  12'd390,  -12'd75,  12'd159,  12'd250,  -12'd242,  12'd159,  12'd232,  12'd588,  -12'd130,  12'd68,  
12'd191,  12'd111,  12'd260,  -12'd115,  -12'd152,  12'd258,  12'd335,  12'd176,  12'd104,  12'd56,  12'd154,  12'd221,  12'd346,  12'd174,  -12'd207,  12'd338,  
12'd2,  12'd103,  -12'd40,  12'd19,  -12'd92,  12'd38,  12'd165,  12'd205,  12'd206,  -12'd1,  -12'd92,  12'd144,  12'd93,  -12'd112,  12'd163,  12'd93,  
-12'd168,  -12'd77,  12'd20,  -12'd14,  12'd202,  -12'd140,  -12'd183,  -12'd32,  -12'd343,  -12'd245,  -12'd56,  -12'd326,  -12'd127,  -12'd324,  -12'd166,  -12'd193,  
-12'd279,  12'd563,  12'd168,  12'd0,  -12'd77,  12'd213,  12'd34,  12'd22,  -12'd315,  -12'd309,  12'd47,  12'd314,  -12'd141,  12'd421,  12'd89,  12'd511,  
-12'd183,  12'd172,  12'd112,  -12'd238,  12'd213,  12'd37,  -12'd128,  -12'd20,  12'd125,  12'd214,  -12'd201,  12'd15,  12'd434,  12'd238,  -12'd339,  -12'd68,  
12'd213,  -12'd124,  -12'd32,  -12'd52,  12'd332,  12'd32,  -12'd262,  -12'd110,  -12'd356,  12'd118,  -12'd109,  12'd64,  -12'd31,  12'd237,  -12'd46,  -12'd109,  
-12'd328,  12'd22,  12'd11,  -12'd89,  12'd60,  -12'd190,  -12'd139,  12'd88,  12'd77,  -12'd170,  12'd239,  12'd128,  -12'd187,  12'd274,  -12'd85,  12'd94,  
-12'd346,  -12'd156,  12'd120,  -12'd171,  -12'd6,  -12'd113,  -12'd33,  12'd372,  12'd181,  12'd122,  12'd69,  -12'd337,  -12'd99,  -12'd300,  12'd198,  -12'd106,  
-12'd254,  12'd146,  12'd58,  -12'd93,  12'd78,  12'd9,  -12'd166,  12'd6,  12'd136,  12'd527,  12'd98,  12'd200,  12'd104,  -12'd158,  12'd170,  12'd349,  
12'd20,  12'd118,  -12'd338,  -12'd160,  12'd172,  12'd233,  12'd240,  12'd161,  -12'd279,  12'd263,  -12'd187,  12'd238,  -12'd467,  -12'd245,  12'd170,  12'd86,  
-12'd58,  12'd44,  12'd360,  -12'd45,  12'd166,  12'd86,  -12'd330,  -12'd331,  12'd31,  12'd188,  12'd57,  12'd334,  -12'd89,  -12'd162,  -12'd383,  12'd104,  
-12'd371,  12'd449,  12'd20,  12'd137,  12'd327,  12'd50,  12'd37,  12'd279,  12'd21,  12'd377,  12'd264,  12'd22,  -12'd130,  -12'd253,  -12'd198,  12'd90,  
-12'd361,  12'd145,  -12'd95,  -12'd26,  12'd10,  12'd209,  -12'd309,  -12'd0,  12'd84,  12'd248,  -12'd23,  -12'd131,  -12'd83,  -12'd180,  -12'd106,  12'd24,  
12'd103,  -12'd238,  -12'd21,  12'd231,  12'd103,  12'd22,  12'd22,  -12'd5,  12'd320,  -12'd128,  12'd57,  12'd0,  -12'd185,  12'd118,  -12'd312,  12'd419,  
12'd282,  12'd228,  12'd30,  12'd65,  -12'd167,  12'd223,  12'd316,  12'd320,  12'd116,  -12'd194,  12'd221,  12'd282,  12'd280,  12'd416,  12'd177,  12'd336,  
12'd163,  12'd238,  12'd147,  12'd27,  12'd84,  12'd236,  12'd133,  -12'd404,  12'd173,  12'd381,  -12'd60,  12'd113,  -12'd75,  12'd30,  12'd208,  12'd104,  
-12'd90,  12'd214,  -12'd370,  12'd88,  12'd132,  12'd157,  12'd48,  12'd0,  -12'd181,  -12'd76,  -12'd116,  -12'd48,  -12'd343,  -12'd371,  12'd356,  -12'd177,  
-12'd388,  12'd267,  12'd89,  -12'd278,  12'd372,  12'd36,  -12'd18,  12'd62,  12'd108,  -12'd72,  -12'd181,  12'd352,  -12'd264,  12'd124,  -12'd38,  -12'd249,  
12'd189,  12'd124,  12'd499,  12'd142,  -12'd66,  12'd410,  -12'd11,  12'd61,  12'd134,  12'd82,  12'd184,  12'd51,  12'd63,  12'd267,  -12'd20,  -12'd101,  
12'd270,  12'd28,  12'd33,  -12'd27,  -12'd388,  12'd351,  -12'd301,  12'd438,  12'd111,  12'd25,  -12'd168,  -12'd107,  12'd38,  12'd654,  -12'd157,  -12'd53,  
-12'd25,  12'd27,  12'd97,  12'd394,  12'd131,  12'd56,  -12'd268,  12'd290,  -12'd189,  12'd66,  -12'd76,  -12'd65,  12'd241,  12'd18,  12'd250,  12'd7,  
12'd163,  -12'd176,  -12'd257,  12'd181,  12'd117,  12'd294,  12'd68,  12'd62,  -12'd158,  -12'd340,  12'd347,  12'd123,  12'd500,  -12'd578,  12'd58,  -12'd0,  
12'd271,  12'd40,  -12'd57,  -12'd184,  -12'd46,  -12'd145,  12'd193,  12'd160,  12'd320,  -12'd40,  12'd71,  12'd339,  -12'd71,  -12'd67,  -12'd43,  -12'd314,  
12'd274,  -12'd171,  12'd114,  12'd48,  -12'd309,  12'd107,  -12'd218,  -12'd285,  12'd196,  -12'd45,  12'd68,  12'd307,  12'd365,  12'd389,  -12'd442,  12'd219,  

12'd48,  -12'd41,  -12'd297,  12'd264,  12'd150,  -12'd107,  -12'd73,  12'd18,  -12'd228,  12'd337,  12'd165,  -12'd80,  -12'd24,  -12'd208,  12'd35,  12'd220,  
-12'd59,  -12'd423,  -12'd77,  12'd180,  12'd117,  12'd168,  -12'd268,  12'd308,  12'd172,  -12'd29,  -12'd382,  -12'd278,  12'd372,  -12'd228,  12'd93,  12'd15,  
-12'd404,  -12'd69,  12'd234,  -12'd144,  12'd275,  -12'd137,  -12'd11,  12'd180,  -12'd191,  12'd186,  12'd51,  12'd267,  -12'd143,  -12'd220,  12'd21,  -12'd324,  
-12'd418,  -12'd702,  12'd241,  -12'd269,  -12'd86,  -12'd204,  12'd56,  -12'd160,  -12'd123,  -12'd133,  12'd268,  12'd21,  -12'd392,  12'd352,  12'd373,  -12'd303,  
12'd40,  12'd103,  12'd72,  12'd138,  -12'd502,  12'd111,  -12'd40,  12'd146,  12'd50,  -12'd133,  -12'd123,  12'd60,  -12'd409,  12'd37,  12'd358,  -12'd208,  
-12'd108,  12'd183,  -12'd44,  -12'd67,  -12'd27,  -12'd260,  12'd4,  -12'd189,  12'd126,  -12'd510,  12'd213,  12'd122,  12'd293,  -12'd353,  12'd180,  12'd249,  
-12'd113,  12'd546,  12'd133,  12'd159,  12'd328,  -12'd53,  12'd35,  -12'd212,  -12'd314,  -12'd197,  -12'd171,  12'd101,  12'd30,  -12'd409,  12'd174,  12'd445,  
-12'd29,  -12'd158,  -12'd76,  12'd273,  12'd169,  -12'd269,  -12'd127,  12'd104,  12'd144,  12'd111,  -12'd324,  12'd315,  -12'd134,  12'd82,  12'd8,  12'd206,  
12'd110,  -12'd65,  12'd82,  12'd178,  -12'd35,  -12'd12,  -12'd43,  -12'd53,  12'd41,  -12'd82,  12'd321,  12'd194,  12'd12,  -12'd341,  12'd285,  -12'd463,  
12'd544,  12'd211,  12'd242,  -12'd0,  12'd133,  12'd62,  12'd25,  -12'd246,  12'd92,  -12'd22,  -12'd136,  -12'd236,  12'd370,  12'd211,  12'd142,  -12'd48,  
12'd44,  12'd210,  -12'd0,  -12'd224,  -12'd596,  12'd192,  12'd167,  12'd14,  12'd315,  12'd50,  12'd367,  -12'd264,  12'd162,  12'd83,  -12'd290,  -12'd37,  
12'd62,  12'd452,  -12'd30,  -12'd77,  12'd16,  12'd230,  -12'd58,  12'd276,  12'd127,  12'd244,  -12'd411,  12'd450,  12'd88,  12'd114,  -12'd42,  -12'd72,  
-12'd149,  12'd332,  12'd119,  -12'd118,  12'd106,  12'd118,  12'd6,  12'd416,  -12'd123,  12'd186,  -12'd260,  -12'd198,  12'd358,  -12'd77,  12'd143,  -12'd370,  
-12'd708,  -12'd225,  -12'd111,  12'd40,  -12'd98,  12'd91,  -12'd453,  -12'd16,  12'd30,  -12'd109,  -12'd306,  12'd47,  12'd295,  -12'd623,  12'd195,  12'd304,  
-12'd260,  -12'd389,  -12'd304,  -12'd93,  12'd110,  -12'd368,  12'd2,  12'd192,  12'd280,  -12'd75,  -12'd126,  -12'd120,  12'd92,  12'd299,  -12'd110,  -12'd13,  
12'd20,  -12'd225,  12'd418,  12'd363,  -12'd286,  12'd413,  12'd4,  12'd192,  12'd117,  12'd46,  12'd182,  -12'd242,  -12'd142,  12'd36,  12'd96,  -12'd395,  
12'd462,  12'd133,  -12'd207,  -12'd72,  -12'd148,  12'd17,  -12'd50,  12'd57,  -12'd145,  -12'd69,  -12'd68,  12'd156,  -12'd336,  -12'd214,  12'd166,  -12'd145,  
12'd79,  12'd432,  -12'd154,  -12'd98,  -12'd19,  12'd37,  -12'd130,  12'd150,  -12'd196,  -12'd187,  12'd229,  -12'd9,  -12'd214,  -12'd192,  12'd365,  -12'd398,  
-12'd104,  12'd133,  -12'd23,  12'd297,  12'd421,  12'd1,  -12'd207,  -12'd90,  12'd73,  -12'd179,  -12'd78,  12'd401,  -12'd63,  12'd22,  12'd25,  -12'd78,  
-12'd142,  -12'd178,  12'd118,  12'd364,  -12'd259,  -12'd8,  -12'd2,  12'd0,  12'd126,  -12'd222,  -12'd13,  12'd68,  -12'd311,  12'd375,  12'd37,  12'd68,  
-12'd6,  -12'd48,  -12'd240,  -12'd218,  -12'd100,  12'd184,  12'd276,  12'd56,  12'd159,  12'd310,  12'd124,  -12'd9,  12'd86,  12'd78,  -12'd55,  -12'd215,  
12'd241,  12'd167,  -12'd276,  -12'd260,  12'd89,  -12'd66,  -12'd527,  -12'd53,  12'd120,  12'd166,  12'd144,  12'd30,  -12'd250,  -12'd432,  12'd76,  -12'd149,  
12'd100,  -12'd105,  -12'd281,  -12'd1,  12'd15,  12'd209,  -12'd115,  -12'd49,  -12'd8,  -12'd17,  12'd53,  12'd412,  12'd125,  -12'd361,  12'd224,  12'd9,  
12'd428,  -12'd12,  12'd439,  -12'd62,  -12'd209,  12'd40,  -12'd66,  12'd276,  12'd585,  12'd98,  12'd4,  12'd4,  -12'd200,  -12'd101,  -12'd122,  12'd44,  
12'd123,  12'd658,  12'd330,  12'd11,  -12'd251,  -12'd287,  12'd56,  -12'd116,  12'd373,  -12'd633,  -12'd61,  12'd78,  -12'd43,  12'd264,  12'd52,  -12'd150,  

-12'd201,  -12'd97,  12'd42,  12'd22,  12'd107,  12'd101,  12'd207,  12'd84,  -12'd245,  12'd358,  -12'd63,  12'd246,  12'd47,  12'd11,  12'd189,  -12'd226,  
12'd260,  -12'd9,  -12'd308,  12'd360,  12'd595,  12'd570,  -12'd63,  12'd346,  12'd245,  12'd317,  -12'd12,  12'd170,  12'd118,  -12'd246,  -12'd92,  12'd23,  
12'd321,  -12'd90,  -12'd25,  12'd55,  -12'd207,  -12'd83,  12'd327,  12'd287,  -12'd20,  -12'd88,  -12'd284,  12'd162,  12'd227,  -12'd558,  12'd199,  12'd195,  
12'd215,  12'd92,  -12'd44,  -12'd52,  12'd203,  12'd207,  12'd387,  -12'd82,  -12'd358,  -12'd270,  12'd299,  12'd246,  12'd531,  12'd165,  12'd186,  12'd284,  
-12'd148,  12'd153,  12'd35,  -12'd43,  12'd171,  -12'd126,  12'd289,  -12'd77,  12'd74,  12'd271,  -12'd135,  12'd61,  -12'd261,  12'd117,  12'd276,  -12'd248,  
-12'd29,  12'd308,  12'd119,  12'd372,  -12'd102,  -12'd283,  -12'd180,  -12'd152,  -12'd215,  -12'd220,  12'd562,  12'd43,  12'd43,  12'd378,  12'd172,  12'd62,  
12'd175,  12'd416,  -12'd91,  12'd152,  12'd561,  -12'd189,  12'd67,  -12'd362,  12'd149,  -12'd127,  12'd117,  12'd186,  -12'd128,  -12'd662,  -12'd303,  12'd176,  
12'd72,  12'd82,  -12'd100,  -12'd320,  12'd61,  -12'd307,  12'd231,  -12'd199,  12'd605,  12'd206,  12'd221,  12'd325,  -12'd188,  -12'd133,  -12'd188,  12'd578,  
12'd333,  12'd210,  12'd49,  12'd78,  -12'd146,  -12'd196,  12'd48,  -12'd215,  12'd239,  -12'd67,  12'd458,  -12'd203,  12'd235,  -12'd195,  12'd46,  -12'd11,  
-12'd169,  12'd356,  -12'd397,  12'd7,  -12'd354,  12'd220,  12'd14,  -12'd159,  12'd359,  -12'd389,  12'd213,  -12'd515,  12'd24,  12'd451,  12'd74,  12'd128,  
12'd78,  12'd167,  12'd339,  12'd133,  -12'd727,  12'd62,  12'd376,  12'd56,  12'd28,  -12'd171,  12'd237,  -12'd309,  -12'd16,  -12'd82,  -12'd103,  12'd287,  
12'd108,  12'd267,  -12'd333,  -12'd537,  -12'd29,  12'd62,  -12'd76,  -12'd314,  -12'd127,  -12'd210,  -12'd185,  -12'd64,  -12'd488,  12'd273,  -12'd278,  12'd99,  
12'd131,  12'd327,  -12'd50,  -12'd293,  -12'd132,  -12'd135,  -12'd76,  12'd109,  -12'd190,  12'd299,  -12'd150,  -12'd382,  12'd126,  12'd553,  12'd249,  -12'd301,  
-12'd3,  12'd98,  -12'd140,  -12'd83,  12'd414,  -12'd89,  -12'd125,  -12'd95,  -12'd189,  12'd120,  -12'd1,  -12'd38,  -12'd190,  12'd123,  12'd164,  -12'd186,  
-12'd421,  12'd102,  12'd3,  -12'd124,  12'd333,  12'd102,  -12'd107,  12'd153,  -12'd127,  12'd34,  -12'd306,  -12'd274,  -12'd272,  12'd411,  12'd393,  12'd265,  
12'd44,  -12'd511,  12'd14,  -12'd450,  -12'd165,  -12'd6,  12'd109,  -12'd66,  12'd218,  12'd208,  -12'd18,  -12'd300,  -12'd21,  12'd129,  -12'd514,  -12'd416,  
12'd111,  12'd312,  12'd298,  -12'd45,  -12'd432,  -12'd145,  12'd275,  -12'd105,  -12'd332,  12'd32,  -12'd146,  -12'd218,  -12'd105,  12'd144,  12'd108,  -12'd289,  
-12'd213,  -12'd221,  12'd129,  -12'd460,  12'd121,  12'd151,  12'd280,  12'd65,  12'd71,  -12'd103,  12'd146,  12'd89,  -12'd323,  12'd121,  -12'd205,  12'd269,  
-12'd614,  -12'd178,  -12'd589,  12'd248,  12'd378,  12'd267,  12'd20,  -12'd241,  12'd65,  -12'd457,  -12'd315,  -12'd57,  -12'd231,  -12'd124,  12'd238,  -12'd101,  
-12'd135,  12'd134,  12'd238,  -12'd55,  12'd103,  12'd250,  12'd202,  -12'd371,  12'd229,  -12'd183,  -12'd217,  12'd184,  -12'd332,  -12'd121,  12'd267,  -12'd118,  
-12'd358,  -12'd54,  12'd107,  12'd379,  12'd191,  12'd79,  12'd409,  12'd237,  12'd343,  12'd139,  -12'd313,  -12'd110,  12'd208,  12'd125,  12'd358,  -12'd192,  
12'd164,  12'd49,  12'd90,  12'd49,  -12'd102,  -12'd156,  -12'd358,  12'd42,  -12'd100,  12'd271,  -12'd244,  12'd203,  -12'd380,  -12'd445,  12'd16,  -12'd145,  
-12'd26,  -12'd103,  -12'd0,  -12'd271,  -12'd92,  12'd90,  -12'd213,  -12'd26,  -12'd127,  12'd445,  -12'd212,  12'd168,  -12'd237,  -12'd206,  -12'd133,  12'd133,  
12'd185,  12'd272,  12'd273,  -12'd211,  -12'd158,  12'd127,  -12'd95,  -12'd106,  12'd90,  12'd172,  -12'd359,  12'd39,  -12'd21,  12'd154,  -12'd78,  -12'd229,  
12'd668,  12'd267,  12'd777,  12'd474,  -12'd442,  12'd514,  12'd13,  -12'd16,  12'd491,  -12'd301,  -12'd169,  12'd160,  12'd298,  -12'd20,  -12'd266,  -12'd239,  

12'd19,  -12'd232,  -12'd312,  12'd6,  -12'd172,  12'd56,  -12'd76,  -12'd31,  12'd221,  -12'd209,  12'd136,  -12'd27,  -12'd101,  -12'd75,  -12'd62,  -12'd111,  
-12'd322,  12'd274,  12'd31,  -12'd487,  12'd45,  -12'd305,  12'd131,  -12'd192,  12'd183,  12'd6,  12'd16,  -12'd254,  12'd60,  -12'd8,  -12'd204,  12'd100,  
12'd138,  12'd13,  -12'd39,  -12'd199,  12'd113,  -12'd282,  -12'd229,  -12'd34,  -12'd96,  -12'd38,  -12'd95,  -12'd225,  -12'd361,  -12'd54,  -12'd30,  -12'd254,  
12'd199,  -12'd215,  -12'd125,  -12'd255,  -12'd38,  -12'd118,  12'd61,  -12'd145,  -12'd288,  -12'd66,  -12'd371,  12'd66,  -12'd166,  -12'd378,  -12'd49,  12'd36,  
-12'd7,  -12'd260,  12'd15,  12'd286,  -12'd54,  12'd289,  -12'd424,  12'd283,  -12'd189,  12'd182,  12'd90,  -12'd59,  -12'd251,  12'd101,  -12'd26,  12'd62,  
12'd168,  -12'd221,  12'd179,  12'd222,  -12'd345,  12'd46,  12'd196,  -12'd205,  -12'd382,  -12'd219,  12'd111,  -12'd151,  -12'd131,  12'd135,  12'd20,  12'd127,  
-12'd58,  -12'd217,  -12'd38,  -12'd26,  -12'd344,  -12'd69,  -12'd85,  -12'd26,  -12'd62,  -12'd237,  -12'd122,  -12'd253,  12'd88,  12'd213,  12'd93,  -12'd175,  
-12'd387,  -12'd12,  -12'd183,  -12'd171,  -12'd200,  -12'd60,  -12'd150,  -12'd227,  -12'd261,  -12'd254,  -12'd147,  12'd189,  12'd69,  -12'd77,  -12'd421,  12'd148,  
-12'd163,  -12'd55,  -12'd93,  12'd49,  12'd198,  -12'd167,  -12'd73,  -12'd116,  -12'd264,  -12'd138,  12'd100,  12'd212,  -12'd47,  -12'd79,  12'd42,  -12'd120,  
12'd30,  -12'd216,  -12'd189,  -12'd229,  -12'd120,  -12'd71,  -12'd191,  12'd81,  12'd79,  -12'd169,  -12'd225,  12'd64,  12'd247,  12'd206,  12'd157,  -12'd114,  
-12'd373,  12'd36,  -12'd7,  -12'd191,  12'd88,  12'd47,  -12'd132,  -12'd76,  12'd70,  -12'd57,  -12'd214,  12'd45,  12'd82,  12'd94,  -12'd127,  -12'd345,  
-12'd87,  -12'd308,  12'd8,  -12'd412,  -12'd289,  12'd84,  12'd172,  -12'd115,  -12'd106,  12'd77,  12'd272,  -12'd9,  12'd135,  12'd79,  -12'd452,  -12'd390,  
12'd80,  -12'd386,  12'd320,  -12'd9,  -12'd273,  -12'd319,  12'd97,  -12'd25,  -12'd261,  12'd201,  -12'd119,  12'd145,  12'd9,  12'd296,  12'd15,  -12'd279,  
12'd349,  12'd43,  12'd11,  -12'd342,  -12'd213,  -12'd94,  -12'd73,  -12'd178,  -12'd22,  12'd150,  12'd165,  -12'd125,  -12'd53,  -12'd199,  12'd127,  12'd52,  
-12'd78,  -12'd2,  12'd62,  12'd204,  -12'd117,  -12'd210,  -12'd291,  -12'd165,  -12'd93,  -12'd17,  -12'd71,  12'd264,  12'd78,  -12'd92,  12'd119,  -12'd58,  
12'd325,  -12'd387,  -12'd230,  12'd96,  -12'd444,  12'd46,  12'd153,  -12'd295,  -12'd66,  -12'd238,  12'd180,  12'd78,  -12'd116,  -12'd191,  -12'd198,  -12'd61,  
12'd58,  12'd115,  12'd92,  12'd183,  -12'd104,  -12'd338,  12'd222,  12'd159,  -12'd104,  12'd60,  -12'd143,  12'd117,  12'd55,  -12'd279,  -12'd42,  -12'd196,  
-12'd144,  -12'd104,  -12'd76,  -12'd293,  -12'd84,  -12'd107,  12'd104,  -12'd67,  -12'd28,  -12'd62,  12'd261,  -12'd277,  -12'd54,  -12'd9,  -12'd211,  12'd116,  
-12'd287,  12'd214,  12'd275,  12'd20,  12'd97,  -12'd180,  -12'd339,  -12'd135,  -12'd239,  -12'd324,  12'd145,  -12'd186,  12'd15,  12'd47,  12'd246,  12'd75,  
-12'd208,  -12'd219,  -12'd250,  -12'd306,  -12'd158,  12'd154,  12'd220,  12'd1,  -12'd327,  12'd80,  12'd146,  12'd281,  -12'd117,  -12'd273,  12'd35,  -12'd62,  
12'd101,  -12'd272,  12'd109,  -12'd173,  -12'd201,  -12'd242,  12'd138,  12'd133,  -12'd63,  -12'd191,  -12'd36,  12'd213,  -12'd24,  -12'd99,  12'd76,  -12'd37,  
-12'd127,  -12'd434,  -12'd17,  12'd6,  -12'd59,  12'd141,  -12'd230,  -12'd388,  -12'd56,  -12'd70,  12'd157,  -12'd175,  12'd28,  12'd20,  -12'd364,  -12'd29,  
-12'd175,  -12'd115,  12'd253,  12'd97,  12'd244,  -12'd94,  -12'd268,  -12'd82,  12'd17,  -12'd111,  12'd299,  -12'd337,  -12'd310,  -12'd4,  12'd66,  -12'd345,  
-12'd116,  -12'd10,  12'd172,  -12'd43,  12'd187,  12'd97,  -12'd162,  12'd44,  -12'd45,  12'd2,  12'd99,  -12'd47,  -12'd268,  -12'd412,  -12'd7,  12'd49,  
-12'd278,  -12'd4,  -12'd82,  -12'd150,  12'd25,  -12'd346,  12'd210,  12'd101,  -12'd322,  12'd16,  -12'd2,  -12'd511,  12'd68,  12'd85,  -12'd125,  12'd49,  

12'd86,  -12'd208,  12'd164,  -12'd421,  -12'd124,  -12'd178,  12'd365,  -12'd14,  12'd16,  -12'd46,  -12'd394,  -12'd50,  -12'd119,  12'd87,  -12'd60,  -12'd68,  
12'd443,  12'd291,  -12'd26,  -12'd379,  -12'd427,  12'd463,  12'd535,  12'd96,  12'd66,  -12'd26,  -12'd46,  -12'd0,  12'd340,  12'd522,  12'd23,  -12'd28,  
12'd70,  -12'd140,  -12'd106,  12'd79,  -12'd77,  12'd129,  12'd413,  -12'd13,  12'd64,  -12'd205,  12'd285,  12'd109,  12'd58,  12'd185,  12'd1,  12'd185,  
12'd237,  12'd246,  12'd108,  12'd68,  12'd487,  12'd593,  -12'd218,  12'd111,  12'd495,  12'd69,  12'd54,  -12'd155,  12'd197,  -12'd92,  12'd244,  -12'd8,  
12'd171,  12'd49,  12'd23,  -12'd308,  12'd12,  -12'd47,  -12'd96,  12'd346,  -12'd356,  12'd33,  12'd316,  12'd98,  12'd468,  -12'd201,  12'd99,  -12'd87,  
-12'd46,  -12'd455,  12'd148,  -12'd281,  -12'd5,  12'd168,  12'd252,  -12'd11,  -12'd189,  -12'd3,  12'd241,  -12'd135,  -12'd358,  12'd0,  12'd40,  12'd23,  
-12'd52,  12'd53,  12'd250,  -12'd358,  12'd301,  12'd27,  12'd197,  12'd125,  -12'd78,  -12'd29,  12'd460,  12'd141,  12'd219,  12'd214,  -12'd124,  -12'd55,  
12'd114,  -12'd45,  12'd472,  -12'd23,  -12'd113,  12'd312,  12'd118,  12'd182,  12'd156,  -12'd82,  -12'd7,  -12'd425,  -12'd118,  -12'd46,  12'd114,  -12'd244,  
12'd263,  12'd274,  -12'd9,  -12'd189,  -12'd10,  12'd240,  -12'd467,  -12'd129,  12'd61,  -12'd61,  12'd145,  -12'd23,  12'd94,  -12'd250,  -12'd372,  12'd282,  
-12'd432,  -12'd242,  12'd558,  12'd156,  -12'd204,  12'd39,  -12'd23,  -12'd183,  -12'd9,  12'd140,  12'd1,  12'd386,  -12'd76,  -12'd122,  12'd297,  12'd459,  
-12'd228,  12'd379,  -12'd70,  -12'd118,  -12'd458,  -12'd424,  12'd138,  12'd10,  -12'd683,  -12'd215,  -12'd302,  12'd1,  -12'd260,  12'd83,  12'd272,  12'd105,  
12'd328,  -12'd327,  12'd44,  -12'd118,  -12'd252,  -12'd323,  -12'd204,  -12'd447,  -12'd189,  -12'd409,  -12'd1,  12'd199,  -12'd364,  12'd179,  -12'd1,  12'd23,  
-12'd78,  -12'd39,  -12'd10,  12'd26,  -12'd113,  -12'd212,  -12'd1,  12'd61,  12'd171,  -12'd242,  -12'd93,  -12'd111,  -12'd298,  -12'd208,  12'd177,  12'd3,  
-12'd525,  12'd196,  -12'd164,  -12'd179,  12'd331,  -12'd186,  12'd283,  -12'd232,  -12'd147,  12'd162,  12'd32,  12'd98,  -12'd170,  -12'd98,  -12'd153,  -12'd195,  
-12'd242,  -12'd80,  12'd228,  -12'd75,  -12'd296,  12'd419,  12'd79,  -12'd20,  -12'd91,  12'd48,  -12'd31,  12'd133,  -12'd908,  -12'd42,  -12'd102,  12'd15,  
12'd148,  12'd187,  12'd362,  -12'd263,  -12'd293,  -12'd102,  12'd175,  12'd87,  -12'd525,  -12'd234,  -12'd436,  12'd21,  12'd1,  12'd322,  -12'd39,  12'd218,  
12'd261,  -12'd4,  12'd555,  -12'd193,  -12'd101,  12'd336,  12'd483,  12'd294,  12'd55,  -12'd396,  -12'd252,  12'd103,  -12'd419,  12'd507,  12'd244,  12'd32,  
12'd57,  -12'd13,  -12'd345,  12'd12,  -12'd27,  -12'd307,  12'd172,  12'd114,  -12'd405,  -12'd190,  -12'd79,  12'd52,  -12'd587,  12'd82,  -12'd187,  -12'd217,  
-12'd399,  -12'd64,  -12'd254,  12'd118,  -12'd149,  -12'd112,  -12'd63,  -12'd180,  -12'd138,  -12'd107,  -12'd320,  12'd148,  12'd201,  12'd350,  12'd81,  -12'd169,  
-12'd50,  -12'd40,  -12'd82,  -12'd312,  12'd101,  12'd135,  12'd260,  -12'd157,  12'd556,  12'd133,  -12'd130,  -12'd246,  -12'd405,  12'd139,  -12'd165,  -12'd537,  
-12'd31,  -12'd262,  12'd132,  -12'd132,  -12'd66,  12'd13,  12'd46,  12'd114,  -12'd430,  12'd343,  -12'd291,  -12'd293,  -12'd61,  12'd506,  -12'd68,  -12'd56,  
-12'd0,  -12'd203,  12'd94,  12'd415,  12'd219,  12'd472,  -12'd258,  12'd55,  -12'd114,  -12'd7,  -12'd46,  -12'd77,  -12'd143,  -12'd261,  12'd389,  12'd76,  
-12'd130,  12'd210,  -12'd276,  12'd292,  -12'd120,  -12'd43,  12'd102,  -12'd64,  12'd143,  12'd81,  -12'd44,  -12'd281,  12'd128,  12'd59,  12'd203,  -12'd376,  
-12'd269,  -12'd175,  -12'd7,  -12'd186,  12'd383,  -12'd443,  12'd66,  -12'd37,  12'd345,  12'd10,  12'd129,  12'd204,  -12'd4,  12'd30,  12'd28,  -12'd47,  
12'd182,  -12'd190,  -12'd235,  12'd280,  -12'd13,  12'd357,  -12'd143,  -12'd199,  12'd242,  12'd439,  -12'd374,  12'd387,  12'd154,  -12'd12,  12'd2,  -12'd110,  

-12'd513,  12'd5,  -12'd174,  -12'd9,  12'd409,  12'd110,  -12'd130,  -12'd44,  12'd58,  -12'd256,  12'd65,  12'd164,  12'd339,  -12'd135,  12'd30,  12'd249,  
12'd3,  12'd184,  -12'd23,  -12'd13,  12'd506,  -12'd185,  12'd108,  12'd9,  12'd304,  -12'd246,  -12'd226,  12'd266,  -12'd21,  12'd181,  -12'd7,  12'd98,  
-12'd42,  12'd412,  12'd31,  -12'd446,  12'd14,  -12'd1,  12'd94,  -12'd41,  -12'd339,  -12'd262,  -12'd300,  -12'd14,  -12'd186,  12'd677,  -12'd4,  12'd233,  
-12'd255,  12'd305,  -12'd101,  12'd97,  12'd65,  12'd126,  12'd434,  -12'd12,  12'd102,  12'd79,  12'd30,  -12'd324,  -12'd149,  12'd796,  12'd33,  12'd186,  
-12'd59,  12'd151,  -12'd127,  -12'd355,  12'd104,  12'd117,  12'd246,  12'd259,  12'd296,  12'd339,  12'd212,  -12'd151,  -12'd350,  12'd303,  12'd211,  -12'd298,  
-12'd164,  12'd59,  12'd124,  12'd6,  12'd91,  -12'd219,  12'd610,  -12'd172,  -12'd146,  -12'd177,  12'd243,  12'd215,  12'd206,  -12'd81,  -12'd366,  12'd225,  
12'd74,  12'd36,  -12'd112,  -12'd31,  12'd65,  -12'd6,  12'd77,  -12'd26,  -12'd82,  12'd276,  -12'd61,  12'd171,  -12'd174,  -12'd51,  -12'd110,  -12'd111,  
12'd66,  -12'd246,  -12'd39,  -12'd401,  -12'd121,  -12'd194,  12'd61,  -12'd122,  -12'd109,  12'd240,  -12'd347,  12'd193,  -12'd188,  -12'd186,  -12'd148,  -12'd400,  
-12'd166,  -12'd344,  12'd455,  12'd214,  -12'd76,  12'd173,  12'd207,  -12'd456,  -12'd214,  12'd149,  12'd356,  12'd55,  12'd89,  12'd0,  -12'd57,  -12'd200,  
12'd215,  12'd363,  12'd161,  12'd88,  -12'd336,  12'd96,  12'd25,  -12'd132,  12'd181,  12'd128,  -12'd5,  12'd104,  12'd121,  -12'd378,  12'd27,  -12'd63,  
12'd237,  12'd217,  12'd54,  -12'd375,  -12'd388,  12'd42,  12'd127,  -12'd199,  -12'd165,  12'd170,  12'd454,  12'd214,  -12'd276,  -12'd136,  -12'd249,  12'd0,  
-12'd90,  12'd231,  -12'd233,  12'd331,  12'd129,  12'd408,  -12'd62,  12'd54,  12'd242,  -12'd268,  -12'd110,  12'd258,  12'd60,  -12'd47,  12'd257,  12'd379,  
-12'd26,  12'd165,  12'd166,  -12'd66,  -12'd126,  12'd77,  12'd10,  -12'd51,  12'd191,  12'd300,  12'd32,  -12'd61,  12'd184,  12'd220,  -12'd48,  12'd55,  
-12'd156,  12'd7,  12'd228,  12'd198,  -12'd248,  -12'd100,  -12'd111,  -12'd426,  12'd17,  12'd156,  12'd61,  12'd29,  12'd115,  12'd111,  -12'd72,  12'd363,  
12'd307,  -12'd210,  12'd60,  12'd321,  -12'd77,  12'd232,  12'd206,  -12'd100,  12'd106,  12'd164,  12'd271,  12'd185,  12'd82,  -12'd178,  -12'd359,  -12'd251,  
12'd308,  12'd231,  -12'd44,  -12'd147,  -12'd518,  12'd175,  12'd186,  -12'd94,  -12'd357,  -12'd376,  12'd36,  12'd517,  12'd279,  12'd145,  12'd162,  12'd406,  
12'd574,  -12'd325,  12'd74,  12'd39,  12'd124,  12'd90,  12'd38,  -12'd37,  12'd210,  12'd170,  12'd50,  12'd81,  -12'd218,  12'd122,  12'd412,  -12'd230,  
12'd132,  12'd46,  -12'd293,  12'd261,  12'd168,  -12'd69,  -12'd101,  12'd165,  12'd112,  12'd91,  12'd6,  12'd249,  12'd394,  -12'd266,  -12'd211,  12'd298,  
12'd108,  12'd121,  -12'd66,  -12'd111,  12'd297,  -12'd334,  -12'd438,  -12'd183,  12'd58,  12'd19,  12'd78,  -12'd304,  12'd139,  -12'd217,  12'd109,  12'd110,  
12'd230,  12'd250,  12'd133,  -12'd92,  12'd109,  12'd21,  -12'd101,  12'd121,  12'd132,  -12'd75,  12'd339,  12'd194,  12'd3,  12'd149,  -12'd205,  12'd336,  
12'd419,  12'd0,  12'd114,  12'd449,  12'd196,  12'd88,  -12'd14,  12'd239,  -12'd175,  12'd420,  -12'd59,  12'd108,  12'd203,  12'd344,  12'd16,  12'd229,  
12'd96,  -12'd96,  12'd147,  -12'd43,  12'd212,  12'd240,  -12'd288,  12'd379,  -12'd633,  -12'd123,  12'd302,  -12'd224,  12'd97,  12'd241,  -12'd232,  12'd11,  
12'd140,  -12'd59,  -12'd120,  12'd127,  -12'd240,  12'd364,  12'd184,  12'd319,  -12'd534,  -12'd78,  -12'd69,  -12'd84,  12'd89,  -12'd483,  12'd140,  12'd188,  
12'd91,  -12'd35,  -12'd144,  -12'd76,  12'd303,  -12'd320,  -12'd81,  12'd136,  -12'd108,  12'd30,  -12'd111,  -12'd301,  12'd333,  -12'd4,  12'd184,  -12'd193,  
12'd75,  -12'd219,  -12'd491,  -12'd18,  12'd247,  12'd206,  12'd155,  12'd162,  -12'd234,  -12'd76,  12'd125,  12'd324,  12'd417,  -12'd183,  -12'd220,  12'd74,  

12'd529,  12'd139,  12'd327,  12'd380,  -12'd113,  12'd237,  12'd577,  12'd389,  -12'd22,  -12'd230,  12'd90,  -12'd142,  12'd79,  12'd540,  -12'd50,  -12'd200,  
-12'd6,  12'd173,  12'd116,  12'd409,  -12'd264,  12'd189,  -12'd70,  -12'd33,  12'd187,  -12'd104,  12'd266,  12'd523,  12'd28,  12'd222,  12'd21,  12'd261,  
-12'd191,  12'd70,  12'd110,  12'd146,  12'd286,  -12'd115,  12'd257,  -12'd27,  12'd354,  12'd541,  12'd402,  12'd61,  12'd140,  12'd243,  -12'd234,  -12'd74,  
-12'd272,  -12'd200,  12'd657,  12'd17,  -12'd202,  -12'd78,  -12'd359,  12'd341,  -12'd52,  12'd326,  -12'd159,  12'd263,  12'd131,  12'd352,  12'd308,  12'd34,  
-12'd214,  -12'd692,  -12'd203,  -12'd162,  -12'd45,  -12'd329,  -12'd314,  -12'd195,  -12'd650,  12'd100,  12'd114,  -12'd75,  -12'd1,  -12'd93,  -12'd227,  -12'd239,  
12'd126,  -12'd89,  12'd361,  12'd242,  -12'd389,  -12'd26,  -12'd201,  -12'd72,  12'd79,  12'd283,  -12'd73,  12'd67,  12'd248,  12'd33,  12'd57,  12'd176,  
-12'd136,  -12'd46,  12'd401,  12'd410,  -12'd282,  12'd175,  12'd150,  12'd229,  -12'd244,  12'd260,  12'd151,  -12'd352,  12'd291,  -12'd143,  12'd29,  12'd105,  
-12'd7,  12'd29,  -12'd342,  12'd305,  -12'd36,  12'd60,  -12'd315,  12'd97,  -12'd318,  -12'd279,  -12'd96,  -12'd144,  12'd448,  12'd108,  12'd301,  12'd153,  
-12'd247,  12'd165,  12'd179,  12'd235,  -12'd512,  12'd79,  -12'd216,  12'd64,  -12'd345,  -12'd105,  -12'd248,  12'd19,  -12'd489,  12'd415,  12'd71,  -12'd182,  
-12'd91,  -12'd441,  12'd285,  -12'd39,  -12'd489,  -12'd14,  -12'd407,  12'd195,  -12'd155,  12'd139,  12'd181,  12'd181,  -12'd508,  12'd355,  -12'd85,  -12'd492,  
12'd175,  12'd22,  -12'd321,  -12'd216,  12'd80,  12'd33,  12'd255,  -12'd37,  -12'd302,  -12'd49,  12'd595,  -12'd327,  12'd185,  12'd82,  12'd75,  -12'd239,  
-12'd233,  12'd162,  -12'd309,  -12'd95,  -12'd328,  -12'd164,  -12'd600,  -12'd68,  12'd62,  12'd74,  -12'd181,  -12'd415,  12'd151,  -12'd45,  12'd230,  -12'd117,  
-12'd301,  12'd258,  -12'd296,  12'd84,  12'd173,  -12'd379,  12'd133,  -12'd306,  12'd115,  -12'd253,  -12'd198,  -12'd121,  -12'd169,  12'd228,  -12'd110,  -12'd104,  
-12'd421,  12'd138,  12'd245,  -12'd138,  -12'd528,  -12'd220,  -12'd110,  -12'd43,  -12'd348,  -12'd221,  12'd601,  12'd145,  -12'd344,  -12'd117,  -12'd145,  -12'd175,  
12'd262,  12'd126,  12'd82,  -12'd38,  12'd104,  -12'd24,  -12'd174,  -12'd345,  -12'd280,  -12'd460,  -12'd57,  -12'd55,  -12'd196,  -12'd248,  12'd20,  -12'd83,  
-12'd34,  12'd33,  -12'd9,  -12'd318,  -12'd219,  -12'd338,  12'd181,  -12'd114,  12'd48,  -12'd44,  12'd12,  12'd24,  12'd112,  -12'd93,  -12'd58,  -12'd67,  
-12'd358,  -12'd158,  12'd301,  12'd67,  -12'd12,  -12'd264,  -12'd51,  -12'd233,  12'd129,  12'd142,  12'd156,  12'd530,  -12'd210,  -12'd189,  12'd223,  12'd253,  
12'd29,  12'd54,  12'd363,  12'd85,  12'd206,  12'd349,  12'd315,  -12'd17,  12'd635,  12'd611,  -12'd477,  -12'd41,  -12'd99,  12'd368,  12'd149,  -12'd510,  
12'd109,  12'd21,  12'd321,  12'd88,  -12'd149,  12'd86,  12'd73,  12'd8,  12'd108,  12'd55,  -12'd295,  12'd133,  -12'd265,  12'd157,  12'd237,  -12'd544,  
12'd361,  -12'd281,  -12'd23,  -12'd31,  -12'd67,  -12'd103,  -12'd289,  -12'd170,  12'd164,  12'd255,  -12'd211,  12'd21,  12'd297,  -12'd89,  12'd184,  -12'd135,  
12'd205,  -12'd75,  12'd28,  12'd350,  -12'd200,  12'd43,  12'd441,  12'd224,  -12'd21,  -12'd327,  -12'd30,  12'd5,  -12'd17,  -12'd195,  -12'd4,  -12'd41,  
-12'd253,  -12'd60,  12'd127,  12'd512,  -12'd203,  12'd528,  12'd67,  -12'd68,  12'd437,  -12'd31,  12'd71,  12'd260,  12'd175,  12'd159,  -12'd220,  12'd51,  
12'd168,  -12'd68,  12'd42,  12'd444,  12'd487,  12'd338,  12'd152,  -12'd81,  -12'd220,  12'd107,  12'd313,  -12'd212,  12'd316,  12'd124,  -12'd13,  12'd81,  
-12'd325,  12'd248,  -12'd481,  12'd333,  12'd90,  12'd66,  -12'd257,  -12'd10,  12'd132,  12'd229,  12'd136,  -12'd152,  12'd228,  -12'd370,  12'd255,  12'd49,  
-12'd370,  -12'd339,  12'd70,  12'd310,  12'd64,  12'd4,  -12'd106,  -12'd123,  -12'd106,  12'd554,  12'd339,  12'd126,  12'd213,  -12'd563,  12'd215,  -12'd77,  

-12'd247,  12'd33,  12'd200,  12'd326,  -12'd233,  -12'd47,  -12'd238,  12'd147,  -12'd139,  12'd142,  -12'd131,  -12'd438,  12'd474,  -12'd157,  12'd313,  12'd53,  
12'd16,  -12'd72,  12'd52,  12'd43,  12'd82,  -12'd321,  -12'd269,  -12'd0,  12'd243,  -12'd6,  12'd12,  12'd319,  -12'd141,  -12'd60,  12'd132,  -12'd22,  
12'd42,  -12'd70,  12'd289,  12'd84,  12'd71,  -12'd153,  -12'd45,  12'd73,  -12'd92,  12'd55,  12'd70,  12'd49,  12'd323,  12'd331,  -12'd101,  -12'd330,  
-12'd8,  12'd13,  -12'd189,  -12'd199,  12'd22,  -12'd147,  12'd16,  -12'd168,  -12'd16,  -12'd174,  -12'd150,  12'd53,  -12'd146,  12'd37,  -12'd107,  -12'd281,  
12'd321,  12'd183,  -12'd96,  12'd22,  -12'd152,  12'd29,  -12'd128,  -12'd134,  -12'd277,  -12'd136,  12'd56,  12'd343,  -12'd239,  12'd24,  -12'd52,  -12'd96,  
-12'd18,  12'd180,  12'd1,  12'd109,  12'd177,  12'd325,  -12'd320,  -12'd152,  12'd66,  12'd72,  -12'd58,  12'd343,  -12'd96,  -12'd146,  12'd182,  -12'd162,  
-12'd103,  -12'd81,  12'd145,  12'd117,  12'd335,  -12'd199,  12'd18,  12'd92,  12'd143,  -12'd161,  -12'd169,  12'd202,  12'd295,  -12'd125,  12'd62,  -12'd77,  
-12'd194,  12'd121,  -12'd202,  12'd318,  -12'd38,  -12'd98,  12'd171,  -12'd393,  12'd96,  -12'd77,  12'd101,  -12'd0,  12'd249,  12'd327,  -12'd59,  12'd144,  
-12'd96,  -12'd105,  -12'd28,  -12'd44,  12'd453,  12'd34,  12'd71,  -12'd30,  12'd469,  -12'd113,  12'd75,  -12'd85,  12'd12,  -12'd77,  -12'd42,  -12'd314,  
12'd711,  12'd81,  -12'd302,  12'd376,  12'd329,  12'd132,  -12'd46,  12'd60,  -12'd16,  12'd338,  -12'd39,  12'd67,  12'd466,  12'd155,  12'd62,  12'd22,  
-12'd283,  12'd122,  -12'd68,  12'd141,  12'd130,  12'd345,  -12'd160,  12'd153,  12'd24,  -12'd242,  12'd23,  -12'd198,  -12'd73,  12'd33,  12'd249,  12'd240,  
-12'd69,  -12'd37,  -12'd12,  12'd101,  12'd53,  -12'd128,  -12'd123,  12'd414,  -12'd331,  12'd161,  -12'd230,  12'd348,  12'd264,  -12'd417,  12'd180,  12'd301,  
-12'd328,  12'd152,  -12'd192,  12'd189,  -12'd214,  12'd185,  12'd392,  -12'd121,  12'd91,  -12'd120,  12'd417,  -12'd80,  12'd543,  12'd29,  -12'd226,  -12'd47,  
-12'd108,  -12'd254,  -12'd175,  12'd411,  -12'd96,  12'd260,  -12'd42,  -12'd56,  12'd302,  -12'd5,  12'd362,  -12'd0,  12'd327,  -12'd150,  -12'd74,  12'd162,  
-12'd467,  -12'd69,  12'd4,  12'd89,  -12'd42,  12'd139,  -12'd403,  12'd178,  12'd141,  -12'd175,  12'd86,  -12'd252,  12'd303,  12'd96,  12'd229,  -12'd151,  
-12'd165,  12'd274,  -12'd167,  -12'd223,  12'd327,  -12'd310,  -12'd445,  -12'd186,  -12'd48,  12'd509,  12'd309,  -12'd272,  -12'd200,  12'd154,  -12'd445,  -12'd146,  
12'd50,  12'd415,  -12'd163,  -12'd112,  -12'd84,  12'd160,  -12'd176,  12'd122,  12'd55,  12'd205,  12'd242,  -12'd315,  12'd189,  -12'd798,  -12'd315,  -12'd101,  
-12'd64,  12'd194,  -12'd429,  -12'd332,  12'd196,  -12'd89,  12'd44,  -12'd224,  12'd164,  -12'd50,  12'd80,  -12'd351,  -12'd104,  -12'd284,  -12'd190,  12'd377,  
-12'd334,  12'd330,  -12'd67,  -12'd213,  12'd462,  -12'd164,  12'd375,  -12'd232,  12'd468,  12'd145,  -12'd4,  12'd265,  -12'd42,  -12'd167,  12'd262,  12'd312,  
-12'd257,  12'd114,  -12'd492,  12'd66,  12'd14,  -12'd35,  12'd178,  12'd289,  -12'd75,  -12'd265,  12'd5,  12'd78,  -12'd263,  -12'd207,  -12'd296,  -12'd175,  
12'd129,  12'd29,  -12'd558,  12'd114,  -12'd39,  -12'd166,  12'd531,  -12'd405,  12'd252,  12'd109,  12'd158,  12'd320,  12'd78,  -12'd119,  -12'd244,  12'd85,  
12'd48,  12'd204,  -12'd275,  -12'd416,  12'd414,  -12'd228,  12'd189,  -12'd282,  12'd198,  12'd192,  -12'd33,  12'd109,  -12'd80,  -12'd324,  -12'd459,  -12'd20,  
12'd251,  12'd420,  12'd65,  -12'd610,  12'd586,  -12'd102,  12'd191,  -12'd308,  -12'd31,  12'd768,  -12'd410,  -12'd45,  -12'd409,  12'd355,  -12'd299,  12'd157,  
-12'd256,  12'd87,  12'd137,  12'd5,  12'd181,  -12'd154,  12'd471,  -12'd334,  12'd43,  -12'd338,  -12'd464,  -12'd80,  -12'd53,  12'd229,  12'd5,  -12'd248,  
12'd16,  -12'd40,  12'd443,  -12'd190,  -12'd216,  12'd135,  12'd135,  -12'd255,  12'd338,  12'd177,  -12'd327,  12'd91,  -12'd248,  12'd164,  12'd17,  -12'd52,  

-12'd671,  -12'd221,  -12'd339,  12'd148,  12'd77,  12'd24,  -12'd400,  12'd168,  12'd158,  -12'd29,  -12'd251,  -12'd112,  12'd101,  -12'd195,  -12'd78,  12'd242,  
12'd82,  -12'd311,  12'd330,  -12'd251,  12'd101,  -12'd216,  12'd12,  12'd101,  -12'd7,  -12'd305,  -12'd338,  -12'd321,  -12'd26,  12'd207,  -12'd217,  -12'd17,  
-12'd354,  -12'd155,  12'd32,  12'd98,  -12'd162,  -12'd224,  -12'd10,  -12'd40,  -12'd345,  12'd22,  -12'd160,  -12'd199,  -12'd95,  12'd811,  12'd48,  -12'd505,  
12'd201,  -12'd261,  12'd392,  -12'd62,  -12'd302,  -12'd112,  -12'd24,  12'd89,  12'd17,  -12'd252,  12'd72,  -12'd31,  -12'd433,  -12'd18,  12'd108,  -12'd526,  
12'd371,  -12'd2,  -12'd110,  12'd351,  -12'd202,  12'd349,  -12'd204,  12'd136,  12'd160,  12'd194,  12'd81,  12'd6,  12'd349,  -12'd286,  12'd161,  12'd310,  
-12'd130,  12'd190,  -12'd119,  12'd265,  12'd213,  -12'd130,  -12'd390,  -12'd302,  -12'd279,  12'd96,  -12'd59,  12'd67,  -12'd145,  12'd109,  12'd4,  -12'd93,  
12'd20,  -12'd266,  -12'd5,  -12'd253,  12'd236,  -12'd55,  12'd73,  12'd55,  -12'd69,  12'd116,  -12'd107,  12'd305,  -12'd491,  12'd137,  12'd82,  12'd11,  
12'd173,  12'd328,  12'd354,  12'd186,  12'd15,  12'd114,  -12'd324,  12'd214,  12'd147,  12'd109,  12'd20,  -12'd121,  -12'd10,  12'd470,  12'd128,  -12'd238,  
12'd3,  12'd54,  -12'd66,  12'd233,  -12'd289,  12'd314,  -12'd301,  12'd396,  -12'd258,  -12'd84,  -12'd2,  -12'd286,  12'd241,  -12'd22,  12'd23,  -12'd267,  
12'd380,  12'd131,  -12'd191,  12'd160,  12'd4,  12'd190,  -12'd334,  -12'd121,  -12'd127,  12'd586,  12'd180,  -12'd248,  12'd358,  -12'd289,  12'd194,  12'd309,  
12'd45,  -12'd120,  12'd47,  12'd200,  -12'd448,  12'd269,  -12'd520,  12'd219,  12'd202,  12'd6,  12'd343,  12'd199,  12'd132,  -12'd91,  12'd53,  -12'd35,  
12'd122,  -12'd443,  12'd70,  12'd142,  12'd289,  12'd88,  12'd11,  12'd104,  12'd357,  12'd17,  12'd238,  12'd278,  12'd171,  -12'd130,  12'd223,  12'd31,  
-12'd173,  12'd147,  12'd415,  12'd50,  -12'd168,  -12'd212,  12'd55,  -12'd112,  12'd259,  12'd36,  12'd132,  12'd441,  12'd18,  12'd452,  12'd55,  -12'd119,  
-12'd399,  -12'd15,  12'd288,  12'd57,  -12'd100,  12'd0,  12'd271,  -12'd30,  -12'd147,  12'd316,  12'd368,  12'd75,  -12'd62,  -12'd141,  12'd52,  -12'd392,  
-12'd419,  -12'd225,  12'd65,  12'd432,  12'd44,  12'd20,  -12'd345,  -12'd200,  12'd2,  12'd100,  12'd13,  -12'd42,  -12'd125,  -12'd219,  12'd102,  -12'd72,  
12'd221,  12'd133,  12'd102,  -12'd54,  -12'd48,  12'd65,  12'd257,  12'd100,  12'd249,  12'd114,  12'd764,  -12'd286,  12'd451,  -12'd52,  12'd60,  -12'd16,  
-12'd138,  12'd153,  12'd11,  12'd256,  -12'd172,  12'd156,  12'd314,  12'd247,  -12'd22,  12'd79,  12'd3,  12'd246,  -12'd33,  -12'd51,  12'd51,  -12'd246,  
12'd72,  -12'd88,  12'd31,  -12'd94,  -12'd120,  12'd110,  -12'd285,  12'd3,  12'd326,  -12'd119,  12'd199,  -12'd221,  12'd180,  12'd713,  12'd87,  -12'd37,  
-12'd297,  -12'd108,  12'd215,  -12'd23,  12'd89,  -12'd314,  12'd40,  12'd119,  12'd70,  -12'd186,  12'd195,  -12'd165,  12'd93,  12'd87,  12'd241,  12'd281,  
12'd209,  12'd297,  12'd629,  12'd123,  -12'd162,  12'd260,  -12'd0,  -12'd1,  -12'd0,  12'd28,  12'd63,  12'd517,  -12'd39,  -12'd17,  12'd62,  12'd107,  
12'd20,  12'd134,  -12'd309,  -12'd159,  -12'd196,  -12'd251,  12'd777,  -12'd228,  12'd168,  -12'd419,  12'd247,  -12'd151,  -12'd65,  -12'd58,  12'd51,  12'd214,  
12'd185,  12'd37,  12'd73,  -12'd136,  12'd93,  12'd191,  12'd441,  12'd9,  12'd177,  12'd201,  -12'd59,  12'd192,  -12'd90,  12'd230,  -12'd134,  -12'd224,  
-12'd14,  -12'd102,  -12'd271,  -12'd296,  12'd172,  12'd12,  -12'd125,  12'd151,  -12'd46,  -12'd274,  12'd109,  12'd28,  -12'd212,  12'd454,  -12'd124,  12'd326,  
-12'd659,  -12'd53,  12'd187,  -12'd63,  -12'd160,  12'd10,  12'd134,  12'd214,  12'd172,  12'd42,  -12'd371,  12'd259,  -12'd58,  12'd24,  12'd403,  12'd157,  
12'd655,  12'd511,  12'd409,  -12'd329,  12'd27,  12'd55,  -12'd266,  -12'd86,  -12'd157,  -12'd28,  12'd333,  12'd111,  12'd120,  -12'd98,  -12'd88,  12'd310,  

12'd1,  12'd283,  -12'd367,  12'd222,  -12'd211,  12'd299,  -12'd415,  -12'd161,  -12'd4,  12'd190,  12'd434,  12'd66,  12'd460,  -12'd197,  -12'd22,  -12'd251,  
12'd118,  -12'd141,  12'd4,  12'd123,  12'd102,  12'd363,  -12'd149,  -12'd367,  12'd155,  12'd56,  -12'd70,  12'd126,  12'd290,  -12'd485,  -12'd254,  -12'd53,  
12'd255,  -12'd145,  -12'd168,  -12'd85,  12'd314,  12'd332,  12'd161,  -12'd299,  -12'd303,  -12'd200,  12'd207,  12'd50,  12'd323,  -12'd130,  -12'd381,  -12'd260,  
12'd253,  12'd452,  12'd111,  12'd217,  12'd288,  12'd141,  -12'd125,  12'd80,  12'd244,  -12'd48,  12'd157,  -12'd86,  -12'd329,  12'd348,  12'd153,  12'd191,  
-12'd103,  12'd80,  12'd210,  12'd27,  -12'd383,  -12'd30,  -12'd106,  -12'd91,  -12'd69,  -12'd2,  -12'd182,  -12'd198,  -12'd681,  -12'd465,  12'd339,  -12'd178,  
12'd113,  12'd142,  -12'd606,  12'd29,  -12'd190,  12'd25,  12'd170,  12'd124,  12'd237,  -12'd183,  12'd395,  12'd129,  12'd188,  -12'd306,  -12'd356,  -12'd19,  
12'd51,  12'd147,  -12'd271,  12'd143,  -12'd235,  -12'd126,  12'd117,  12'd153,  -12'd69,  12'd10,  12'd260,  12'd290,  12'd418,  -12'd368,  -12'd566,  12'd167,  
12'd295,  12'd428,  -12'd101,  -12'd251,  -12'd28,  -12'd73,  12'd297,  -12'd433,  12'd199,  -12'd273,  12'd81,  12'd81,  12'd224,  12'd409,  -12'd124,  12'd459,  
-12'd28,  12'd366,  12'd319,  -12'd421,  12'd281,  12'd202,  12'd125,  12'd55,  -12'd56,  12'd62,  -12'd120,  -12'd207,  -12'd67,  12'd541,  -12'd266,  -12'd173,  
12'd82,  12'd235,  12'd238,  12'd123,  -12'd297,  12'd75,  12'd287,  12'd293,  -12'd236,  -12'd3,  12'd105,  -12'd188,  -12'd526,  -12'd59,  12'd31,  -12'd560,  
-12'd154,  -12'd353,  -12'd237,  -12'd471,  -12'd86,  -12'd474,  12'd232,  -12'd108,  -12'd135,  -12'd129,  12'd332,  -12'd146,  -12'd293,  -12'd180,  12'd201,  -12'd217,  
-12'd81,  -12'd416,  -12'd229,  12'd80,  -12'd395,  -12'd81,  -12'd301,  -12'd318,  12'd78,  12'd5,  12'd210,  12'd18,  -12'd187,  12'd89,  -12'd616,  12'd224,  
-12'd2,  -12'd90,  -12'd352,  -12'd431,  12'd353,  -12'd246,  12'd178,  -12'd245,  12'd184,  12'd436,  12'd32,  -12'd161,  12'd127,  12'd222,  -12'd169,  -12'd172,  
12'd30,  12'd143,  12'd242,  -12'd419,  12'd130,  -12'd209,  12'd145,  -12'd323,  12'd203,  12'd31,  12'd56,  -12'd81,  12'd8,  12'd523,  -12'd258,  -12'd145,  
12'd615,  12'd301,  -12'd25,  12'd178,  -12'd180,  -12'd5,  12'd286,  12'd162,  12'd235,  12'd123,  12'd274,  -12'd171,  -12'd81,  -12'd253,  -12'd32,  -12'd97,  
-12'd172,  -12'd111,  12'd84,  12'd178,  -12'd244,  -12'd111,  -12'd43,  -12'd291,  -12'd38,  -12'd166,  -12'd59,  12'd108,  -12'd288,  -12'd104,  -12'd10,  -12'd322,  
12'd106,  -12'd438,  -12'd291,  -12'd346,  12'd166,  -12'd250,  -12'd292,  -12'd315,  12'd250,  -12'd180,  12'd116,  12'd182,  12'd60,  -12'd97,  -12'd255,  -12'd299,  
-12'd18,  -12'd270,  12'd30,  -12'd150,  12'd73,  -12'd481,  12'd120,  -12'd254,  12'd305,  12'd69,  -12'd246,  12'd380,  -12'd221,  -12'd170,  -12'd122,  -12'd173,  
12'd90,  -12'd251,  12'd114,  -12'd9,  12'd112,  -12'd51,  -12'd208,  12'd58,  12'd418,  12'd73,  -12'd296,  -12'd244,  12'd76,  12'd451,  12'd19,  -12'd327,  
12'd33,  -12'd66,  -12'd506,  -12'd236,  -12'd110,  12'd318,  -12'd47,  12'd265,  12'd606,  12'd272,  12'd84,  12'd194,  12'd184,  -12'd484,  12'd408,  -12'd227,  
12'd253,  12'd0,  12'd198,  12'd211,  -12'd495,  12'd103,  -12'd54,  -12'd78,  12'd12,  -12'd497,  12'd158,  12'd52,  12'd130,  -12'd91,  -12'd27,  12'd23,  
12'd124,  -12'd341,  -12'd371,  12'd371,  -12'd373,  12'd228,  -12'd109,  12'd97,  12'd16,  -12'd26,  12'd338,  12'd4,  12'd91,  -12'd24,  -12'd69,  12'd333,  
12'd197,  12'd90,  12'd4,  12'd234,  -12'd288,  12'd396,  12'd41,  12'd92,  12'd77,  -12'd188,  12'd409,  -12'd72,  12'd433,  12'd65,  12'd200,  -12'd19,  
-12'd358,  12'd121,  12'd224,  12'd170,  12'd383,  12'd268,  -12'd260,  -12'd71,  -12'd46,  12'd500,  12'd142,  -12'd100,  12'd151,  -12'd480,  12'd147,  12'd266,  
-12'd333,  -12'd194,  12'd125,  12'd146,  -12'd30,  12'd328,  12'd49,  12'd128,  12'd147,  12'd408,  12'd374,  12'd320,  12'd196,  -12'd123,  12'd80,  12'd153,  

-12'd270,  -12'd277,  12'd70,  12'd218,  -12'd25,  12'd84,  -12'd55,  -12'd234,  12'd69,  12'd75,  12'd69,  -12'd30,  -12'd297,  -12'd117,  12'd279,  12'd48,  
12'd32,  12'd109,  12'd102,  -12'd138,  12'd72,  -12'd300,  12'd98,  -12'd137,  -12'd115,  -12'd130,  -12'd2,  -12'd330,  12'd97,  12'd166,  -12'd7,  -12'd188,  
12'd198,  -12'd108,  -12'd284,  12'd78,  12'd168,  -12'd433,  -12'd11,  12'd9,  -12'd35,  -12'd102,  -12'd104,  12'd68,  12'd159,  12'd279,  12'd46,  -12'd140,  
12'd194,  -12'd82,  -12'd136,  12'd192,  -12'd243,  12'd259,  -12'd215,  12'd22,  -12'd73,  12'd109,  -12'd174,  -12'd119,  -12'd254,  12'd264,  12'd145,  -12'd269,  
12'd239,  12'd10,  12'd31,  -12'd201,  -12'd23,  -12'd55,  12'd7,  12'd370,  12'd122,  -12'd290,  -12'd184,  12'd94,  12'd1,  12'd150,  -12'd55,  -12'd316,  
12'd8,  -12'd20,  12'd319,  -12'd253,  -12'd182,  12'd367,  -12'd15,  -12'd114,  -12'd139,  12'd257,  -12'd213,  12'd142,  12'd88,  -12'd291,  -12'd109,  -12'd68,  
12'd184,  12'd204,  -12'd62,  -12'd107,  -12'd62,  -12'd244,  -12'd195,  -12'd143,  12'd335,  -12'd337,  -12'd119,  -12'd256,  -12'd182,  -12'd439,  12'd307,  -12'd417,  
12'd65,  12'd78,  -12'd52,  -12'd198,  -12'd193,  -12'd102,  -12'd65,  12'd4,  -12'd52,  -12'd238,  12'd227,  12'd193,  12'd198,  -12'd61,  12'd106,  12'd145,  
12'd162,  12'd241,  12'd93,  -12'd142,  -12'd37,  12'd27,  -12'd378,  12'd202,  -12'd209,  -12'd211,  12'd103,  -12'd426,  12'd104,  -12'd92,  -12'd183,  -12'd419,  
-12'd64,  -12'd75,  12'd51,  12'd67,  -12'd188,  12'd71,  -12'd46,  -12'd29,  -12'd280,  -12'd162,  -12'd225,  12'd247,  12'd76,  -12'd155,  12'd145,  -12'd281,  
12'd193,  12'd68,  12'd104,  12'd115,  12'd74,  12'd74,  -12'd148,  12'd2,  -12'd53,  -12'd149,  -12'd60,  12'd21,  12'd55,  -12'd195,  -12'd96,  12'd15,  
12'd191,  -12'd143,  12'd192,  12'd369,  -12'd145,  12'd28,  -12'd324,  -12'd314,  12'd69,  -12'd60,  -12'd87,  -12'd304,  12'd347,  -12'd13,  -12'd72,  -12'd113,  
12'd108,  12'd89,  -12'd171,  -12'd197,  12'd45,  -12'd368,  12'd191,  -12'd290,  12'd272,  12'd282,  12'd211,  -12'd193,  -12'd77,  -12'd139,  -12'd379,  -12'd84,  
12'd51,  -12'd237,  12'd102,  12'd232,  -12'd153,  -12'd114,  -12'd40,  12'd132,  12'd317,  -12'd190,  12'd69,  -12'd231,  12'd109,  12'd189,  12'd343,  12'd136,  
12'd165,  -12'd314,  12'd42,  12'd63,  -12'd114,  12'd13,  12'd198,  12'd133,  -12'd77,  -12'd159,  -12'd54,  -12'd88,  -12'd207,  12'd166,  12'd27,  -12'd142,  
-12'd74,  12'd25,  12'd286,  -12'd121,  -12'd139,  -12'd240,  12'd54,  -12'd10,  12'd20,  12'd101,  -12'd105,  -12'd128,  -12'd132,  -12'd137,  -12'd24,  -12'd141,  
12'd124,  -12'd74,  -12'd164,  -12'd268,  12'd89,  -12'd250,  -12'd67,  12'd80,  -12'd192,  12'd138,  -12'd105,  12'd101,  -12'd301,  12'd219,  -12'd71,  -12'd58,  
-12'd47,  -12'd170,  -12'd29,  -12'd28,  -12'd10,  12'd53,  -12'd208,  -12'd233,  12'd45,  -12'd191,  -12'd8,  -12'd232,  12'd0,  -12'd55,  -12'd244,  12'd77,  
12'd125,  -12'd69,  -12'd145,  -12'd181,  -12'd314,  12'd198,  -12'd2,  -12'd113,  -12'd39,  12'd17,  12'd76,  -12'd294,  -12'd80,  -12'd444,  -12'd41,  -12'd56,  
12'd387,  -12'd234,  -12'd135,  -12'd129,  -12'd130,  -12'd28,  -12'd28,  -12'd70,  12'd124,  -12'd18,  12'd14,  12'd43,  12'd261,  12'd187,  -12'd15,  -12'd411,  
12'd88,  -12'd22,  -12'd38,  -12'd354,  -12'd97,  12'd315,  -12'd22,  -12'd57,  -12'd5,  12'd280,  -12'd305,  -12'd65,  -12'd216,  12'd130,  12'd167,  -12'd92,  
-12'd69,  -12'd435,  -12'd258,  -12'd22,  -12'd164,  -12'd107,  -12'd110,  12'd221,  12'd164,  -12'd9,  -12'd254,  -12'd178,  -12'd330,  -12'd371,  -12'd1,  12'd228,  
-12'd120,  -12'd72,  12'd147,  12'd29,  12'd76,  12'd150,  -12'd88,  -12'd291,  12'd44,  -12'd120,  -12'd268,  -12'd415,  -12'd206,  12'd258,  -12'd226,  12'd5,  
12'd125,  12'd121,  -12'd155,  -12'd298,  12'd321,  -12'd299,  -12'd158,  -12'd207,  12'd210,  12'd270,  -12'd180,  12'd37,  -12'd106,  -12'd69,  -12'd198,  -12'd22,  
12'd151,  12'd27,  -12'd47,  -12'd21,  -12'd86,  -12'd54,  -12'd199,  -12'd241,  -12'd51,  12'd77,  -12'd30,  -12'd100,  -12'd194,  12'd250,  -12'd244,  -12'd47,  

12'd130,  -12'd37,  -12'd383,  -12'd302,  -12'd230,  -12'd643,  12'd635,  -12'd495,  12'd53,  -12'd577,  -12'd503,  -12'd38,  -12'd299,  12'd226,  -12'd466,  -12'd413,  
-12'd35,  12'd211,  -12'd431,  -12'd78,  -12'd88,  -12'd362,  -12'd7,  12'd13,  12'd13,  12'd267,  -12'd520,  -12'd41,  -12'd379,  -12'd260,  -12'd70,  -12'd423,  
12'd405,  12'd254,  -12'd389,  -12'd28,  -12'd80,  12'd399,  -12'd500,  12'd293,  -12'd61,  12'd77,  12'd82,  12'd134,  12'd38,  -12'd759,  12'd277,  12'd238,  
12'd49,  -12'd181,  -12'd92,  12'd106,  12'd143,  12'd114,  -12'd2,  -12'd76,  12'd234,  12'd170,  12'd200,  12'd283,  12'd56,  -12'd390,  12'd175,  12'd79,  
-12'd583,  12'd237,  12'd27,  -12'd187,  -12'd40,  12'd106,  12'd1,  -12'd214,  -12'd70,  -12'd139,  12'd182,  12'd100,  -12'd213,  12'd60,  12'd91,  12'd258,  
-12'd87,  -12'd10,  -12'd317,  12'd20,  -12'd379,  -12'd95,  12'd7,  12'd45,  -12'd210,  12'd148,  -12'd217,  -12'd15,  12'd63,  -12'd47,  -12'd221,  -12'd402,  
12'd330,  12'd150,  12'd160,  -12'd155,  12'd115,  -12'd46,  -12'd54,  12'd229,  12'd63,  -12'd95,  -12'd329,  -12'd148,  -12'd234,  -12'd30,  12'd124,  -12'd18,  
12'd117,  -12'd82,  -12'd40,  -12'd209,  -12'd333,  -12'd107,  12'd21,  12'd442,  12'd112,  12'd34,  -12'd73,  12'd57,  -12'd234,  -12'd670,  12'd449,  -12'd127,  
12'd257,  -12'd250,  12'd20,  12'd43,  -12'd62,  12'd161,  12'd69,  12'd33,  -12'd61,  -12'd176,  -12'd223,  -12'd259,  12'd86,  12'd165,  -12'd37,  12'd47,  
-12'd436,  -12'd132,  -12'd177,  12'd138,  -12'd127,  12'd75,  12'd358,  12'd204,  12'd308,  -12'd315,  12'd409,  12'd175,  -12'd21,  12'd336,  -12'd105,  -12'd156,  
12'd308,  12'd157,  12'd370,  -12'd24,  12'd295,  -12'd37,  12'd47,  -12'd125,  -12'd114,  -12'd5,  -12'd738,  12'd95,  -12'd84,  12'd348,  12'd76,  12'd61,  
-12'd21,  -12'd164,  12'd398,  -12'd113,  12'd227,  12'd101,  -12'd350,  12'd161,  12'd3,  12'd44,  -12'd422,  12'd133,  12'd91,  12'd179,  12'd16,  -12'd420,  
12'd56,  -12'd42,  12'd353,  12'd212,  -12'd132,  -12'd1,  12'd140,  -12'd212,  12'd16,  -12'd164,  12'd181,  -12'd76,  -12'd249,  -12'd177,  12'd91,  12'd59,  
12'd169,  12'd285,  12'd99,  -12'd384,  12'd93,  -12'd217,  -12'd61,  -12'd79,  12'd173,  12'd71,  12'd237,  -12'd304,  -12'd53,  12'd334,  -12'd236,  12'd126,  
-12'd113,  12'd1,  12'd191,  -12'd183,  12'd9,  12'd78,  12'd11,  12'd215,  12'd113,  -12'd434,  12'd195,  -12'd134,  12'd79,  12'd541,  12'd356,  -12'd35,  
12'd30,  12'd12,  12'd224,  12'd130,  -12'd117,  -12'd41,  -12'd586,  12'd58,  -12'd365,  12'd97,  -12'd437,  12'd18,  12'd17,  12'd179,  -12'd54,  -12'd3,  
-12'd73,  -12'd22,  12'd261,  12'd169,  -12'd23,  -12'd46,  12'd16,  -12'd45,  -12'd81,  -12'd140,  -12'd245,  12'd50,  -12'd32,  12'd128,  -12'd3,  -12'd194,  
-12'd147,  12'd575,  12'd283,  -12'd414,  12'd303,  -12'd213,  12'd131,  -12'd123,  -12'd152,  12'd127,  -12'd8,  12'd136,  -12'd84,  -12'd38,  12'd356,  -12'd91,  
-12'd40,  12'd45,  12'd324,  -12'd4,  -12'd50,  -12'd118,  12'd258,  -12'd362,  12'd69,  -12'd335,  -12'd322,  12'd325,  12'd63,  12'd304,  -12'd417,  -12'd44,  
12'd176,  12'd340,  -12'd186,  -12'd294,  -12'd317,  -12'd8,  -12'd146,  12'd154,  -12'd186,  -12'd484,  -12'd228,  -12'd261,  12'd73,  12'd216,  -12'd484,  -12'd583,  
-12'd334,  12'd37,  12'd208,  12'd217,  12'd505,  12'd178,  -12'd282,  12'd18,  -12'd152,  12'd102,  12'd199,  -12'd1,  -12'd71,  -12'd18,  -12'd65,  -12'd162,  
12'd71,  12'd28,  -12'd48,  -12'd261,  12'd52,  -12'd110,  -12'd387,  -12'd104,  -12'd179,  -12'd377,  12'd148,  12'd127,  12'd128,  -12'd100,  12'd15,  12'd229,  
12'd400,  -12'd361,  -12'd90,  12'd288,  -12'd74,  -12'd50,  -12'd171,  -12'd167,  12'd367,  12'd135,  -12'd90,  12'd164,  -12'd16,  -12'd283,  -12'd80,  12'd9,  
12'd457,  -12'd103,  12'd252,  12'd121,  -12'd104,  -12'd147,  12'd96,  12'd171,  12'd150,  12'd191,  12'd24,  12'd397,  12'd90,  12'd154,  -12'd345,  12'd41,  
12'd93,  -12'd238,  -12'd359,  -12'd261,  -12'd263,  -12'd327,  -12'd73,  12'd230,  12'd467,  -12'd526,  -12'd266,  -12'd510,  12'd25,  12'd207,  -12'd100,  -12'd71,  

12'd61,  -12'd137,  -12'd53,  12'd6,  12'd17,  12'd261,  -12'd579,  12'd8,  12'd112,  -12'd45,  12'd197,  -12'd258,  -12'd47,  -12'd524,  12'd29,  -12'd122,  
-12'd28,  12'd132,  -12'd78,  12'd221,  12'd6,  -12'd139,  -12'd151,  -12'd27,  12'd464,  12'd138,  -12'd279,  -12'd415,  12'd193,  -12'd85,  -12'd96,  12'd637,  
-12'd68,  -12'd283,  -12'd68,  -12'd353,  12'd383,  12'd34,  -12'd51,  12'd352,  12'd52,  12'd27,  -12'd463,  12'd150,  12'd152,  -12'd1,  -12'd82,  12'd143,  
-12'd361,  -12'd458,  -12'd216,  -12'd166,  12'd223,  -12'd221,  12'd69,  -12'd83,  -12'd56,  -12'd475,  -12'd195,  -12'd233,  -12'd163,  12'd577,  -12'd274,  12'd158,  
-12'd174,  -12'd73,  12'd190,  -12'd212,  12'd218,  -12'd6,  -12'd199,  12'd27,  -12'd75,  -12'd70,  -12'd225,  12'd332,  -12'd333,  12'd168,  12'd106,  -12'd473,  
12'd79,  12'd134,  -12'd302,  -12'd161,  12'd433,  -12'd278,  -12'd190,  12'd247,  -12'd28,  -12'd265,  -12'd47,  -12'd37,  12'd24,  -12'd573,  12'd168,  -12'd100,  
-12'd45,  12'd12,  -12'd42,  -12'd382,  12'd31,  -12'd129,  12'd170,  -12'd15,  -12'd1,  12'd231,  -12'd207,  12'd248,  -12'd190,  12'd51,  12'd187,  12'd110,  
12'd411,  -12'd203,  12'd179,  -12'd115,  12'd163,  12'd102,  12'd128,  12'd340,  -12'd35,  12'd349,  -12'd62,  12'd466,  -12'd188,  12'd354,  12'd278,  12'd223,  
12'd603,  -12'd341,  12'd362,  12'd126,  12'd5,  12'd286,  12'd105,  12'd315,  -12'd30,  -12'd143,  12'd89,  12'd283,  -12'd52,  12'd489,  12'd147,  12'd275,  
12'd441,  12'd284,  -12'd93,  12'd8,  12'd289,  12'd226,  -12'd52,  -12'd108,  12'd26,  -12'd457,  -12'd383,  -12'd289,  12'd290,  12'd348,  -12'd120,  -12'd75,  
-12'd39,  -12'd68,  -12'd14,  12'd117,  12'd132,  12'd183,  -12'd122,  12'd158,  12'd295,  -12'd17,  12'd43,  -12'd313,  12'd98,  -12'd258,  12'd170,  12'd100,  
12'd115,  -12'd213,  -12'd224,  -12'd157,  -12'd274,  12'd176,  -12'd91,  12'd243,  12'd268,  12'd159,  12'd5,  12'd54,  12'd451,  12'd225,  -12'd10,  -12'd5,  
-12'd16,  -12'd156,  -12'd440,  12'd443,  -12'd272,  -12'd135,  -12'd26,  12'd104,  -12'd47,  12'd245,  12'd378,  12'd286,  12'd195,  -12'd356,  12'd123,  12'd339,  
-12'd34,  -12'd562,  12'd449,  12'd184,  12'd119,  12'd84,  12'd114,  12'd406,  -12'd195,  12'd0,  12'd144,  12'd254,  12'd405,  -12'd394,  12'd86,  -12'd23,  
-12'd62,  -12'd193,  -12'd286,  -12'd82,  -12'd262,  -12'd92,  12'd316,  12'd346,  -12'd83,  12'd109,  -12'd20,  -12'd310,  12'd413,  -12'd45,  -12'd27,  12'd361,  
-12'd51,  -12'd257,  12'd338,  -12'd35,  12'd292,  -12'd17,  -12'd348,  12'd146,  12'd52,  -12'd12,  -12'd7,  -12'd5,  12'd149,  -12'd230,  -12'd22,  -12'd168,  
-12'd251,  12'd73,  12'd25,  12'd75,  12'd119,  -12'd179,  -12'd262,  12'd155,  12'd165,  -12'd127,  -12'd186,  12'd148,  12'd118,  12'd42,  -12'd4,  12'd270,  
-12'd153,  -12'd177,  -12'd258,  12'd41,  -12'd11,  -12'd201,  12'd6,  -12'd229,  -12'd244,  -12'd65,  -12'd77,  12'd56,  -12'd271,  -12'd224,  -12'd184,  12'd36,  
12'd250,  12'd339,  12'd102,  -12'd179,  -12'd528,  12'd331,  -12'd210,  12'd13,  12'd123,  12'd125,  12'd236,  12'd99,  -12'd100,  -12'd58,  12'd105,  12'd85,  
-12'd169,  12'd67,  -12'd131,  -12'd9,  12'd378,  -12'd154,  12'd91,  12'd365,  12'd123,  -12'd262,  12'd52,  12'd247,  -12'd105,  12'd135,  12'd218,  -12'd74,  
-12'd64,  12'd81,  -12'd155,  12'd322,  12'd183,  12'd173,  -12'd147,  -12'd140,  -12'd26,  -12'd157,  -12'd63,  12'd378,  12'd87,  12'd80,  -12'd137,  -12'd154,  
12'd91,  12'd115,  -12'd362,  12'd65,  -12'd279,  -12'd222,  -12'd442,  -12'd305,  12'd82,  12'd194,  12'd119,  -12'd6,  -12'd206,  12'd118,  12'd145,  12'd126,  
-12'd17,  -12'd145,  -12'd86,  -12'd405,  12'd149,  -12'd254,  12'd224,  12'd222,  12'd161,  12'd268,  -12'd187,  12'd132,  -12'd200,  12'd303,  12'd160,  -12'd96,  
12'd85,  -12'd233,  12'd479,  -12'd146,  12'd85,  12'd84,  12'd264,  -12'd137,  12'd428,  -12'd181,  -12'd109,  12'd215,  -12'd202,  12'd78,  12'd150,  12'd41,  
12'd25,  -12'd95,  12'd201,  -12'd114,  12'd96,  -12'd154,  12'd393,  12'd312,  -12'd208,  -12'd618,  -12'd56,  12'd247,  12'd46,  -12'd5,  -12'd121,  12'd129,  

12'd387,  12'd175,  -12'd299,  -12'd143,  -12'd177,  12'd436,  -12'd202,  12'd119,  -12'd76,  12'd22,  12'd143,  12'd126,  12'd74,  -12'd379,  12'd318,  12'd122,  
-12'd142,  12'd139,  -12'd232,  -12'd205,  -12'd172,  12'd165,  12'd161,  12'd444,  -12'd41,  12'd184,  12'd155,  12'd22,  -12'd69,  -12'd312,  12'd338,  12'd146,  
12'd49,  12'd317,  -12'd368,  12'd114,  12'd160,  12'd122,  -12'd26,  -12'd287,  -12'd169,  12'd42,  12'd26,  12'd83,  -12'd310,  12'd466,  12'd83,  12'd179,  
12'd9,  12'd65,  12'd155,  -12'd346,  -12'd79,  12'd111,  12'd108,  -12'd318,  12'd121,  12'd224,  -12'd204,  -12'd61,  -12'd16,  12'd239,  -12'd151,  -12'd203,  
-12'd125,  -12'd39,  -12'd362,  -12'd65,  12'd390,  12'd80,  -12'd175,  -12'd328,  -12'd382,  -12'd280,  -12'd55,  -12'd114,  -12'd433,  12'd265,  12'd208,  12'd277,  
12'd239,  -12'd168,  -12'd28,  12'd152,  12'd26,  -12'd220,  12'd178,  12'd161,  -12'd131,  12'd362,  12'd25,  -12'd15,  12'd168,  -12'd95,  -12'd90,  12'd284,  
12'd138,  12'd264,  -12'd74,  12'd178,  12'd207,  -12'd9,  12'd165,  -12'd333,  -12'd6,  12'd371,  -12'd325,  -12'd241,  12'd30,  12'd56,  -12'd55,  12'd384,  
-12'd73,  12'd21,  -12'd184,  -12'd148,  12'd14,  -12'd307,  -12'd303,  12'd167,  -12'd304,  12'd172,  12'd324,  12'd179,  12'd211,  -12'd196,  12'd32,  12'd270,  
12'd226,  -12'd332,  12'd62,  12'd88,  -12'd92,  -12'd105,  -12'd170,  -12'd279,  12'd49,  -12'd116,  -12'd70,  12'd42,  -12'd160,  12'd108,  -12'd291,  12'd279,  
12'd487,  12'd530,  12'd105,  -12'd253,  -12'd41,  12'd96,  12'd146,  -12'd86,  12'd105,  -12'd148,  -12'd96,  12'd394,  12'd224,  -12'd195,  -12'd358,  -12'd324,  
-12'd239,  12'd312,  -12'd134,  -12'd104,  12'd109,  -12'd65,  -12'd100,  12'd111,  12'd42,  12'd324,  12'd224,  12'd20,  12'd40,  -12'd28,  -12'd272,  -12'd52,  
12'd283,  12'd233,  12'd210,  -12'd18,  -12'd58,  12'd200,  -12'd235,  12'd181,  12'd118,  12'd92,  -12'd28,  12'd18,  -12'd60,  -12'd149,  -12'd75,  12'd214,  
12'd352,  12'd190,  12'd156,  12'd58,  -12'd171,  12'd438,  12'd167,  12'd72,  12'd323,  -12'd52,  12'd286,  12'd170,  -12'd177,  -12'd359,  -12'd94,  12'd38,  
12'd307,  -12'd514,  12'd76,  -12'd51,  12'd176,  12'd105,  12'd85,  -12'd138,  12'd313,  12'd228,  12'd36,  -12'd116,  -12'd100,  12'd76,  12'd356,  12'd158,  
12'd152,  12'd61,  -12'd451,  12'd270,  -12'd28,  12'd223,  -12'd10,  -12'd141,  12'd89,  12'd281,  12'd17,  -12'd38,  12'd193,  -12'd61,  -12'd32,  12'd237,  
12'd123,  -12'd51,  -12'd107,  -12'd105,  -12'd264,  12'd49,  -12'd87,  -12'd253,  12'd271,  -12'd177,  -12'd435,  12'd98,  12'd73,  12'd262,  12'd60,  -12'd231,  
12'd312,  12'd174,  12'd201,  12'd331,  12'd63,  12'd117,  12'd27,  -12'd118,  12'd203,  12'd7,  -12'd56,  -12'd39,  12'd100,  12'd429,  12'd52,  -12'd23,  
-12'd288,  12'd118,  -12'd101,  12'd196,  -12'd201,  12'd90,  12'd45,  -12'd269,  12'd430,  12'd196,  -12'd77,  -12'd87,  12'd77,  -12'd551,  -12'd96,  12'd43,  
-12'd187,  -12'd117,  12'd42,  12'd47,  12'd33,  12'd177,  12'd108,  12'd103,  -12'd188,  12'd100,  12'd334,  -12'd171,  12'd94,  -12'd363,  12'd104,  -12'd337,  
-12'd433,  -12'd0,  -12'd160,  12'd121,  12'd89,  12'd49,  -12'd122,  -12'd140,  -12'd91,  12'd126,  12'd89,  12'd134,  12'd133,  12'd6,  -12'd29,  12'd104,  
12'd278,  -12'd71,  12'd405,  12'd232,  -12'd212,  12'd206,  -12'd8,  12'd354,  -12'd9,  12'd18,  -12'd348,  12'd202,  12'd100,  12'd375,  12'd155,  12'd10,  
12'd216,  12'd212,  12'd56,  12'd144,  12'd214,  -12'd180,  -12'd407,  12'd535,  -12'd50,  -12'd185,  -12'd250,  -12'd14,  12'd335,  12'd281,  12'd35,  12'd3,  
-12'd441,  -12'd146,  12'd22,  12'd141,  12'd264,  12'd111,  12'd87,  12'd11,  -12'd557,  -12'd872,  12'd88,  12'd73,  12'd208,  -12'd347,  12'd95,  -12'd188,  
-12'd349,  12'd122,  -12'd365,  -12'd88,  -12'd219,  -12'd2,  -12'd91,  12'd87,  12'd192,  -12'd401,  12'd28,  12'd204,  -12'd94,  -12'd10,  12'd256,  -12'd260,  
-12'd170,  12'd179,  12'd119,  12'd197,  -12'd92,  -12'd53,  12'd162,  -12'd49,  12'd11,  -12'd260,  12'd177,  12'd270,  12'd116,  -12'd94,  -12'd62,  12'd19,  

12'd226,  12'd199,  12'd84,  12'd149,  -12'd534,  12'd168,  12'd613,  -12'd14,  12'd92,  -12'd260,  -12'd389,  12'd288,  -12'd485,  12'd46,  -12'd225,  12'd44,  
12'd59,  12'd40,  -12'd217,  -12'd352,  -12'd217,  12'd163,  -12'd233,  -12'd265,  12'd189,  12'd65,  12'd502,  -12'd80,  -12'd315,  12'd300,  -12'd260,  -12'd156,  
12'd105,  12'd66,  -12'd543,  -12'd140,  12'd217,  12'd77,  -12'd236,  -12'd240,  -12'd174,  12'd190,  12'd94,  -12'd200,  -12'd211,  12'd278,  -12'd215,  12'd269,  
-12'd187,  12'd179,  12'd3,  12'd192,  12'd246,  -12'd91,  -12'd152,  -12'd108,  12'd120,  12'd124,  -12'd31,  -12'd57,  12'd46,  12'd25,  -12'd79,  -12'd108,  
12'd172,  12'd615,  12'd170,  -12'd173,  12'd99,  12'd217,  -12'd91,  12'd266,  -12'd168,  12'd64,  12'd96,  12'd160,  12'd298,  12'd94,  12'd201,  12'd268,  
12'd118,  -12'd80,  12'd113,  -12'd45,  12'd32,  12'd212,  -12'd126,  -12'd11,  -12'd101,  12'd158,  -12'd246,  12'd185,  -12'd30,  12'd689,  -12'd136,  12'd133,  
12'd192,  -12'd77,  12'd140,  12'd154,  -12'd281,  12'd41,  -12'd77,  12'd246,  12'd65,  12'd92,  -12'd209,  -12'd335,  12'd396,  12'd344,  12'd415,  -12'd19,  
-12'd472,  -12'd268,  12'd54,  -12'd356,  -12'd149,  -12'd228,  -12'd130,  -12'd42,  12'd214,  12'd18,  12'd260,  -12'd1,  -12'd225,  -12'd116,  12'd59,  -12'd149,  
-12'd503,  -12'd189,  -12'd55,  -12'd214,  -12'd105,  12'd391,  -12'd303,  12'd185,  -12'd4,  -12'd31,  -12'd139,  12'd251,  -12'd47,  -12'd70,  12'd145,  -12'd174,  
-12'd138,  12'd286,  -12'd241,  -12'd54,  12'd178,  12'd120,  12'd140,  12'd97,  12'd217,  12'd232,  -12'd208,  -12'd219,  -12'd156,  12'd73,  -12'd62,  12'd47,  
12'd223,  12'd105,  -12'd67,  12'd446,  12'd102,  12'd683,  -12'd570,  12'd342,  -12'd373,  12'd245,  -12'd217,  12'd255,  12'd227,  12'd149,  12'd224,  12'd244,  
-12'd198,  12'd509,  12'd145,  12'd228,  12'd270,  -12'd159,  -12'd468,  12'd321,  12'd22,  -12'd253,  12'd523,  12'd347,  -12'd201,  12'd93,  12'd14,  12'd410,  
-12'd234,  -12'd157,  12'd122,  12'd221,  12'd35,  12'd175,  -12'd178,  12'd389,  12'd364,  -12'd614,  12'd131,  -12'd81,  12'd95,  -12'd4,  12'd66,  -12'd16,  
-12'd83,  12'd9,  -12'd326,  12'd40,  -12'd376,  12'd4,  -12'd48,  -12'd15,  12'd161,  12'd20,  12'd8,  12'd88,  12'd60,  -12'd44,  -12'd290,  12'd213,  
12'd85,  12'd20,  -12'd312,  -12'd19,  12'd42,  12'd26,  -12'd389,  12'd83,  -12'd201,  12'd47,  -12'd26,  -12'd57,  12'd114,  12'd27,  12'd22,  12'd195,  
12'd363,  12'd292,  -12'd72,  -12'd57,  12'd381,  -12'd54,  -12'd362,  12'd263,  -12'd138,  -12'd56,  -12'd298,  12'd259,  12'd200,  12'd282,  -12'd18,  12'd238,  
12'd74,  12'd420,  12'd384,  -12'd136,  12'd291,  12'd331,  12'd168,  -12'd160,  -12'd179,  12'd156,  -12'd22,  -12'd80,  -12'd374,  12'd114,  12'd46,  12'd183,  
12'd35,  12'd94,  12'd46,  -12'd22,  12'd85,  12'd54,  12'd211,  -12'd152,  12'd539,  -12'd16,  -12'd162,  -12'd85,  -12'd257,  -12'd230,  -12'd150,  12'd187,  
-12'd351,  12'd296,  -12'd186,  -12'd155,  12'd221,  -12'd129,  12'd77,  12'd102,  -12'd173,  12'd88,  12'd24,  -12'd40,  -12'd301,  12'd181,  -12'd104,  -12'd134,  
-12'd163,  -12'd298,  12'd221,  -12'd74,  12'd100,  -12'd88,  12'd0,  -12'd232,  -12'd416,  -12'd6,  12'd195,  12'd45,  -12'd214,  12'd12,  -12'd124,  -12'd1,  
12'd404,  -12'd76,  12'd42,  12'd58,  -12'd15,  -12'd183,  12'd153,  12'd152,  12'd300,  -12'd210,  -12'd258,  12'd21,  12'd101,  12'd29,  12'd28,  -12'd36,  
-12'd273,  -12'd154,  12'd0,  12'd23,  12'd16,  -12'd119,  -12'd313,  12'd89,  -12'd68,  12'd207,  -12'd2,  -12'd206,  -12'd88,  -12'd10,  -12'd54,  -12'd5,  
-12'd149,  -12'd136,  12'd156,  12'd58,  -12'd182,  -12'd154,  -12'd332,  12'd101,  -12'd53,  12'd102,  -12'd216,  -12'd45,  -12'd89,  -12'd140,  12'd173,  12'd105,  
-12'd310,  12'd128,  -12'd67,  12'd361,  -12'd59,  12'd198,  -12'd71,  -12'd75,  -12'd91,  -12'd216,  12'd7,  12'd246,  -12'd17,  12'd396,  12'd51,  -12'd119,  
-12'd203,  -12'd241,  -12'd65,  12'd233,  -12'd194,  -12'd183,  -12'd1,  -12'd77,  12'd40,  -12'd417,  -12'd208,  12'd147,  12'd87,  -12'd106,  12'd57,  12'd368,  

-12'd85,  12'd18,  12'd8,  -12'd27,  12'd148,  -12'd87,  -12'd387,  12'd290,  -12'd23,  12'd94,  -12'd484,  -12'd220,  12'd248,  -12'd6,  -12'd399,  -12'd29,  
-12'd333,  12'd133,  12'd365,  12'd168,  12'd355,  -12'd16,  -12'd435,  -12'd225,  -12'd96,  12'd258,  -12'd281,  12'd134,  12'd149,  12'd338,  12'd304,  12'd374,  
12'd35,  -12'd265,  12'd128,  -12'd217,  12'd33,  -12'd218,  -12'd38,  12'd57,  12'd19,  -12'd151,  12'd35,  12'd323,  -12'd123,  12'd391,  12'd274,  12'd317,  
12'd29,  -12'd113,  12'd273,  12'd143,  -12'd9,  12'd103,  12'd204,  12'd195,  -12'd58,  -12'd69,  12'd38,  12'd251,  -12'd223,  12'd522,  12'd326,  -12'd61,  
12'd307,  -12'd232,  12'd15,  -12'd111,  -12'd211,  -12'd168,  12'd308,  -12'd172,  12'd251,  -12'd9,  -12'd60,  12'd134,  -12'd211,  12'd114,  12'd150,  -12'd168,  
-12'd126,  -12'd225,  12'd112,  -12'd28,  12'd133,  12'd122,  -12'd384,  12'd258,  -12'd384,  12'd76,  -12'd264,  -12'd69,  -12'd111,  12'd212,  12'd59,  -12'd297,  
12'd214,  12'd216,  12'd190,  12'd374,  -12'd43,  12'd219,  12'd94,  -12'd73,  12'd118,  12'd4,  12'd221,  12'd428,  -12'd177,  12'd1,  12'd180,  -12'd327,  
-12'd98,  12'd248,  12'd333,  12'd176,  12'd85,  12'd115,  12'd159,  12'd356,  12'd268,  12'd23,  12'd49,  -12'd108,  12'd14,  12'd528,  12'd211,  -12'd357,  
-12'd215,  12'd151,  12'd118,  12'd86,  -12'd135,  12'd79,  12'd118,  12'd155,  -12'd88,  -12'd486,  12'd258,  12'd198,  -12'd368,  12'd40,  12'd128,  -12'd27,  
12'd182,  12'd230,  12'd11,  -12'd242,  12'd184,  12'd71,  12'd140,  -12'd169,  12'd208,  -12'd331,  -12'd27,  -12'd166,  12'd31,  -12'd413,  12'd146,  12'd221,  
12'd321,  12'd2,  -12'd94,  -12'd94,  12'd71,  -12'd242,  -12'd65,  -12'd88,  12'd360,  12'd64,  12'd636,  -12'd170,  -12'd185,  12'd248,  12'd57,  -12'd24,  
12'd32,  12'd270,  12'd89,  -12'd151,  -12'd263,  12'd192,  12'd48,  12'd366,  -12'd166,  12'd74,  12'd149,  -12'd27,  12'd63,  12'd29,  12'd55,  12'd318,  
12'd100,  12'd214,  12'd162,  12'd149,  12'd89,  -12'd89,  12'd66,  12'd223,  -12'd151,  12'd48,  12'd5,  12'd196,  12'd91,  12'd353,  -12'd50,  -12'd125,  
-12'd271,  12'd71,  12'd241,  -12'd12,  -12'd5,  12'd20,  12'd317,  12'd19,  -12'd106,  -12'd113,  12'd342,  12'd92,  -12'd171,  -12'd173,  -12'd119,  -12'd464,  
12'd167,  12'd4,  -12'd125,  12'd149,  12'd154,  12'd95,  12'd117,  12'd51,  -12'd18,  -12'd708,  -12'd215,  -12'd326,  -12'd137,  12'd25,  12'd119,  -12'd341,  
-12'd37,  12'd213,  -12'd85,  -12'd99,  12'd576,  -12'd252,  -12'd359,  12'd27,  12'd309,  -12'd194,  12'd100,  -12'd73,  12'd83,  12'd24,  -12'd427,  12'd38,  
-12'd112,  -12'd315,  -12'd71,  12'd143,  -12'd13,  -12'd18,  12'd268,  -12'd78,  -12'd106,  -12'd97,  12'd142,  12'd107,  -12'd11,  12'd125,  -12'd218,  12'd175,  
12'd289,  -12'd85,  -12'd26,  12'd68,  -12'd116,  12'd449,  -12'd57,  -12'd296,  12'd110,  12'd15,  12'd95,  -12'd304,  12'd173,  12'd202,  12'd100,  -12'd61,  
-12'd13,  -12'd243,  -12'd12,  12'd87,  12'd231,  -12'd409,  -12'd257,  -12'd1,  12'd529,  12'd66,  12'd135,  -12'd130,  -12'd238,  12'd30,  12'd3,  12'd258,  
12'd288,  -12'd54,  12'd81,  -12'd199,  -12'd156,  -12'd168,  -12'd189,  -12'd21,  -12'd9,  12'd127,  -12'd235,  12'd83,  12'd117,  -12'd144,  -12'd132,  -12'd27,  
-12'd290,  -12'd175,  -12'd433,  -12'd73,  -12'd204,  12'd19,  -12'd25,  12'd79,  12'd204,  -12'd191,  12'd508,  -12'd8,  -12'd105,  12'd78,  12'd35,  12'd91,  
-12'd44,  12'd165,  -12'd338,  12'd4,  -12'd125,  12'd190,  12'd216,  -12'd510,  12'd389,  -12'd298,  12'd140,  12'd417,  -12'd310,  12'd105,  12'd8,  12'd116,  
-12'd64,  12'd250,  12'd98,  -12'd376,  -12'd16,  -12'd18,  12'd266,  -12'd177,  12'd213,  12'd307,  12'd113,  -12'd15,  12'd57,  12'd426,  12'd53,  12'd368,  
12'd141,  -12'd12,  12'd335,  12'd276,  -12'd71,  -12'd235,  -12'd110,  -12'd104,  -12'd240,  12'd137,  -12'd258,  -12'd176,  -12'd390,  12'd123,  12'd188,  -12'd127,  
12'd415,  12'd370,  12'd402,  -12'd106,  12'd312,  12'd351,  -12'd228,  12'd86,  -12'd53,  12'd576,  -12'd244,  12'd215,  -12'd91,  12'd247,  12'd109,  12'd89,  

12'd307,  -12'd24,  12'd114,  12'd126,  12'd279,  -12'd81,  12'd184,  12'd96,  12'd158,  12'd36,  -12'd130,  -12'd50,  12'd169,  -12'd241,  12'd95,  12'd125,  
-12'd187,  -12'd82,  12'd127,  -12'd119,  -12'd249,  -12'd93,  12'd599,  12'd196,  12'd65,  -12'd235,  12'd255,  -12'd237,  -12'd71,  12'd142,  -12'd381,  -12'd129,  
-12'd21,  12'd273,  -12'd77,  12'd122,  12'd115,  -12'd4,  -12'd57,  12'd200,  12'd31,  -12'd129,  12'd25,  -12'd179,  -12'd245,  -12'd357,  -12'd52,  -12'd138,  
12'd302,  12'd330,  12'd146,  12'd219,  -12'd142,  -12'd241,  -12'd139,  -12'd85,  -12'd4,  12'd81,  12'd99,  12'd199,  12'd509,  -12'd521,  -12'd2,  -12'd259,  
12'd361,  12'd406,  -12'd277,  12'd241,  -12'd110,  -12'd16,  -12'd28,  -12'd75,  -12'd179,  12'd348,  -12'd222,  12'd131,  12'd204,  12'd170,  -12'd236,  12'd110,  
-12'd166,  -12'd166,  12'd159,  -12'd312,  -12'd104,  -12'd287,  -12'd60,  -12'd32,  12'd226,  -12'd73,  12'd399,  -12'd57,  12'd155,  -12'd61,  12'd113,  -12'd249,  
-12'd138,  -12'd368,  12'd87,  12'd284,  12'd59,  -12'd195,  12'd171,  12'd224,  12'd199,  -12'd302,  12'd176,  12'd342,  12'd101,  12'd341,  12'd181,  -12'd390,  
12'd94,  -12'd279,  12'd117,  12'd221,  -12'd244,  -12'd247,  -12'd301,  12'd41,  12'd279,  -12'd294,  12'd411,  -12'd299,  12'd117,  -12'd44,  12'd78,  12'd71,  
-12'd449,  12'd143,  -12'd419,  12'd124,  12'd167,  -12'd290,  -12'd278,  12'd317,  12'd123,  12'd575,  12'd151,  12'd55,  12'd376,  -12'd398,  12'd204,  12'd268,  
-12'd144,  -12'd225,  -12'd53,  12'd211,  12'd242,  12'd186,  -12'd354,  -12'd53,  -12'd397,  12'd817,  12'd238,  -12'd24,  -12'd48,  -12'd234,  12'd99,  12'd223,  
-12'd112,  12'd82,  -12'd87,  12'd142,  -12'd530,  12'd51,  12'd99,  -12'd168,  -12'd59,  -12'd181,  -12'd374,  -12'd386,  -12'd174,  12'd375,  12'd4,  12'd94,  
12'd75,  -12'd76,  -12'd224,  12'd46,  -12'd188,  12'd150,  -12'd3,  12'd201,  -12'd96,  12'd17,  -12'd309,  -12'd377,  12'd77,  -12'd37,  12'd54,  12'd259,  
-12'd464,  12'd277,  -12'd377,  12'd89,  12'd136,  -12'd112,  12'd174,  12'd209,  12'd448,  12'd252,  12'd10,  -12'd171,  -12'd196,  -12'd160,  12'd267,  12'd310,  
-12'd502,  12'd87,  -12'd546,  -12'd100,  12'd276,  -12'd12,  -12'd90,  12'd91,  -12'd54,  12'd209,  12'd289,  12'd228,  -12'd207,  -12'd112,  -12'd17,  12'd403,  
-12'd135,  -12'd184,  12'd426,  -12'd13,  12'd245,  12'd290,  12'd332,  12'd268,  12'd373,  12'd192,  12'd55,  12'd493,  -12'd51,  -12'd91,  12'd43,  -12'd113,  
12'd145,  -12'd85,  -12'd52,  12'd51,  -12'd69,  12'd136,  12'd40,  12'd204,  12'd153,  -12'd53,  -12'd252,  -12'd166,  -12'd199,  -12'd49,  -12'd216,  12'd153,  
-12'd248,  -12'd12,  -12'd29,  -12'd68,  -12'd219,  12'd187,  12'd96,  12'd383,  -12'd382,  -12'd31,  12'd108,  12'd144,  -12'd34,  12'd28,  12'd222,  -12'd171,  
12'd8,  -12'd409,  -12'd146,  -12'd47,  12'd239,  12'd66,  12'd24,  12'd177,  -12'd273,  -12'd201,  12'd316,  12'd364,  12'd288,  -12'd32,  12'd4,  12'd2,  
12'd133,  12'd469,  -12'd111,  -12'd31,  12'd44,  12'd475,  -12'd230,  -12'd260,  12'd359,  -12'd290,  12'd97,  -12'd125,  12'd263,  12'd157,  12'd17,  -12'd219,  
-12'd34,  -12'd47,  12'd471,  12'd7,  -12'd78,  12'd59,  12'd149,  12'd0,  -12'd124,  -12'd224,  12'd376,  -12'd205,  -12'd152,  12'd261,  12'd91,  12'd25,  
12'd145,  -12'd183,  -12'd276,  -12'd30,  -12'd127,  12'd358,  -12'd124,  -12'd132,  -12'd67,  12'd109,  -12'd4,  12'd44,  -12'd405,  12'd155,  12'd255,  -12'd8,  
-12'd137,  12'd13,  -12'd190,  12'd217,  -12'd131,  12'd442,  12'd129,  -12'd85,  12'd36,  12'd264,  12'd45,  12'd124,  12'd32,  -12'd513,  -12'd72,  -12'd55,  
12'd269,  12'd85,  -12'd396,  -12'd144,  -12'd36,  12'd141,  12'd321,  -12'd333,  -12'd92,  -12'd49,  12'd443,  -12'd40,  -12'd50,  -12'd385,  12'd114,  12'd50,  
-12'd163,  12'd201,  12'd103,  -12'd243,  12'd120,  -12'd198,  12'd429,  -12'd85,  12'd243,  -12'd124,  -12'd49,  -12'd242,  -12'd202,  12'd373,  12'd59,  -12'd39,  
-12'd144,  -12'd75,  -12'd213,  -12'd310,  -12'd230,  12'd45,  -12'd132,  -12'd116,  12'd398,  12'd29,  -12'd239,  -12'd310,  12'd62,  12'd19,  -12'd536,  12'd20,  

-12'd70,  -12'd143,  12'd33,  12'd106,  -12'd144,  12'd138,  12'd63,  12'd145,  -12'd170,  12'd114,  -12'd402,  -12'd440,  12'd83,  12'd102,  -12'd25,  12'd21,  
-12'd426,  12'd9,  12'd153,  -12'd44,  -12'd7,  -12'd181,  -12'd76,  -12'd112,  -12'd262,  -12'd268,  -12'd262,  -12'd183,  -12'd427,  12'd304,  12'd191,  12'd67,  
-12'd34,  -12'd106,  12'd237,  -12'd11,  -12'd181,  12'd274,  -12'd423,  12'd193,  12'd349,  -12'd270,  12'd308,  12'd160,  12'd20,  12'd509,  12'd88,  -12'd132,  
-12'd186,  12'd448,  12'd390,  -12'd181,  -12'd97,  -12'd74,  12'd166,  12'd261,  12'd131,  -12'd71,  12'd61,  -12'd157,  -12'd24,  -12'd561,  12'd226,  12'd291,  
-12'd266,  -12'd263,  -12'd21,  12'd193,  -12'd110,  -12'd465,  -12'd93,  -12'd208,  12'd187,  12'd52,  -12'd11,  -12'd34,  -12'd215,  12'd50,  12'd233,  -12'd403,  
-12'd13,  12'd103,  -12'd424,  12'd4,  12'd170,  12'd127,  -12'd448,  -12'd372,  -12'd125,  12'd54,  -12'd148,  -12'd55,  -12'd68,  -12'd509,  -12'd224,  -12'd319,  
12'd358,  -12'd171,  12'd90,  12'd424,  -12'd164,  -12'd99,  12'd207,  -12'd37,  -12'd456,  12'd204,  12'd168,  -12'd13,  -12'd72,  -12'd198,  -12'd281,  -12'd190,  
12'd87,  -12'd45,  12'd184,  -12'd335,  -12'd389,  -12'd26,  12'd248,  12'd48,  -12'd107,  12'd430,  12'd66,  12'd242,  12'd154,  -12'd41,  -12'd261,  12'd29,  
-12'd77,  -12'd124,  12'd172,  -12'd100,  -12'd304,  -12'd62,  -12'd31,  12'd195,  -12'd290,  12'd10,  -12'd190,  12'd37,  -12'd32,  -12'd92,  12'd191,  -12'd45,  
-12'd555,  12'd256,  12'd433,  -12'd80,  -12'd247,  -12'd454,  -12'd81,  -12'd126,  -12'd52,  12'd297,  12'd155,  12'd66,  -12'd208,  12'd42,  12'd110,  12'd125,  
-12'd99,  12'd29,  -12'd414,  12'd154,  -12'd40,  -12'd180,  -12'd269,  12'd26,  12'd482,  12'd59,  12'd522,  12'd13,  -12'd104,  -12'd433,  12'd64,  12'd246,  
12'd320,  -12'd301,  -12'd462,  12'd171,  -12'd116,  12'd217,  -12'd111,  12'd152,  12'd182,  12'd451,  12'd128,  12'd347,  12'd276,  -12'd624,  -12'd93,  12'd214,  
12'd451,  -12'd134,  12'd88,  12'd295,  12'd409,  -12'd221,  12'd205,  12'd359,  12'd509,  12'd283,  12'd150,  12'd103,  12'd447,  -12'd182,  12'd37,  12'd47,  
-12'd28,  -12'd317,  -12'd110,  12'd220,  -12'd33,  12'd155,  -12'd23,  -12'd136,  12'd180,  12'd333,  -12'd165,  12'd17,  -12'd232,  12'd626,  -12'd3,  -12'd128,  
12'd822,  12'd327,  12'd515,  12'd107,  -12'd678,  12'd224,  -12'd116,  12'd97,  12'd196,  -12'd79,  -12'd193,  12'd33,  12'd437,  -12'd293,  12'd140,  -12'd112,  
12'd175,  -12'd333,  12'd74,  -12'd1,  12'd0,  -12'd264,  12'd467,  -12'd113,  12'd787,  12'd336,  12'd440,  -12'd90,  12'd96,  12'd199,  12'd122,  12'd183,  
-12'd159,  -12'd109,  -12'd123,  12'd10,  -12'd42,  12'd168,  -12'd4,  12'd165,  12'd124,  -12'd57,  12'd662,  12'd208,  12'd295,  12'd273,  12'd264,  -12'd30,  
-12'd310,  12'd279,  -12'd47,  12'd424,  12'd61,  12'd319,  12'd104,  -12'd164,  -12'd354,  -12'd356,  12'd291,  12'd56,  12'd85,  -12'd29,  12'd325,  12'd114,  
-12'd179,  12'd50,  -12'd321,  -12'd25,  12'd153,  -12'd285,  12'd98,  12'd8,  -12'd173,  12'd220,  -12'd264,  -12'd540,  12'd323,  12'd6,  12'd73,  -12'd295,  
12'd430,  -12'd160,  12'd473,  -12'd305,  12'd357,  -12'd374,  -12'd283,  12'd223,  12'd11,  12'd303,  12'd351,  12'd14,  12'd155,  12'd126,  -12'd314,  -12'd69,  
12'd0,  -12'd109,  -12'd169,  -12'd4,  -12'd99,  12'd132,  12'd260,  12'd146,  -12'd142,  -12'd154,  12'd53,  -12'd486,  12'd353,  12'd111,  12'd14,  12'd120,  
-12'd468,  12'd48,  -12'd380,  12'd15,  -12'd247,  -12'd255,  12'd131,  -12'd276,  -12'd76,  -12'd227,  12'd125,  -12'd345,  12'd252,  12'd128,  12'd63,  12'd175,  
-12'd351,  -12'd142,  -12'd152,  -12'd157,  -12'd203,  -12'd17,  -12'd287,  12'd50,  -12'd456,  -12'd189,  12'd59,  -12'd354,  -12'd445,  12'd125,  -12'd236,  12'd375,  
-12'd333,  12'd84,  -12'd583,  12'd120,  -12'd33,  -12'd32,  -12'd85,  12'd49,  12'd11,  -12'd230,  12'd131,  12'd150,  -12'd215,  -12'd418,  12'd78,  -12'd70,  
-12'd770,  12'd309,  -12'd310,  -12'd62,  -12'd174,  -12'd483,  -12'd153,  -12'd118,  -12'd410,  12'd39,  12'd171,  -12'd78,  -12'd339,  12'd178,  -12'd218,  -12'd160,  

12'd47,  -12'd28,  12'd180,  -12'd25,  12'd169,  -12'd135,  -12'd188,  12'd339,  12'd105,  12'd213,  12'd56,  12'd456,  12'd48,  12'd455,  12'd67,  12'd206,  
12'd82,  -12'd134,  12'd113,  12'd82,  12'd30,  12'd201,  12'd286,  12'd123,  12'd267,  -12'd60,  12'd356,  12'd341,  12'd220,  12'd270,  -12'd9,  12'd6,  
12'd293,  12'd98,  -12'd196,  -12'd292,  -12'd464,  -12'd73,  -12'd117,  12'd48,  12'd169,  12'd8,  -12'd47,  12'd25,  12'd289,  12'd194,  -12'd333,  -12'd306,  
12'd242,  12'd201,  -12'd431,  12'd154,  -12'd153,  12'd23,  12'd191,  12'd127,  -12'd270,  12'd9,  12'd297,  -12'd52,  12'd66,  12'd80,  -12'd161,  12'd313,  
12'd403,  12'd604,  -12'd370,  -12'd197,  12'd320,  12'd167,  12'd128,  -12'd68,  -12'd103,  12'd155,  12'd197,  12'd32,  12'd569,  -12'd23,  12'd32,  12'd83,  
-12'd210,  12'd387,  12'd50,  12'd26,  12'd276,  12'd430,  -12'd127,  -12'd142,  12'd144,  12'd10,  -12'd167,  12'd450,  12'd6,  12'd322,  12'd156,  12'd142,  
12'd69,  12'd24,  12'd116,  12'd412,  12'd99,  -12'd189,  12'd42,  -12'd127,  -12'd171,  12'd11,  12'd368,  12'd131,  12'd56,  -12'd30,  12'd94,  -12'd177,  
-12'd481,  -12'd267,  12'd104,  12'd60,  -12'd177,  12'd183,  12'd196,  -12'd2,  12'd360,  -12'd374,  -12'd13,  -12'd236,  12'd181,  -12'd250,  12'd58,  12'd69,  
-12'd142,  12'd119,  -12'd66,  12'd42,  12'd24,  -12'd309,  -12'd302,  -12'd342,  12'd219,  12'd188,  12'd40,  12'd212,  -12'd56,  -12'd98,  -12'd101,  12'd257,  
12'd13,  -12'd472,  -12'd84,  12'd287,  12'd502,  12'd318,  -12'd35,  12'd54,  -12'd47,  -12'd9,  -12'd237,  -12'd3,  12'd244,  -12'd556,  -12'd239,  12'd408,  
-12'd133,  12'd80,  12'd36,  12'd4,  12'd366,  -12'd50,  12'd105,  -12'd244,  12'd19,  12'd147,  12'd278,  12'd106,  12'd135,  -12'd207,  -12'd54,  12'd343,  
-12'd56,  12'd127,  12'd221,  12'd228,  12'd140,  12'd234,  12'd228,  -12'd30,  -12'd254,  -12'd213,  12'd143,  -12'd63,  -12'd12,  -12'd53,  12'd179,  -12'd168,  
12'd33,  -12'd356,  12'd81,  -12'd181,  -12'd22,  12'd41,  12'd214,  -12'd286,  12'd48,  -12'd162,  -12'd74,  12'd24,  -12'd273,  -12'd131,  -12'd158,  -12'd149,  
-12'd290,  -12'd298,  -12'd482,  12'd99,  -12'd28,  -12'd112,  12'd20,  -12'd260,  12'd199,  -12'd94,  -12'd69,  12'd18,  12'd38,  -12'd29,  12'd240,  -12'd15,  
-12'd184,  -12'd197,  -12'd203,  -12'd20,  12'd135,  12'd64,  -12'd18,  12'd19,  -12'd225,  12'd368,  12'd411,  12'd46,  12'd142,  12'd318,  12'd324,  12'd326,  
12'd18,  12'd164,  12'd10,  -12'd370,  -12'd365,  -12'd76,  12'd220,  -12'd256,  -12'd181,  12'd75,  -12'd222,  12'd59,  -12'd87,  -12'd145,  -12'd130,  12'd272,  
12'd497,  12'd42,  12'd19,  12'd154,  12'd309,  -12'd299,  12'd52,  -12'd225,  -12'd408,  12'd23,  -12'd390,  12'd87,  12'd148,  12'd232,  12'd187,  -12'd30,  
12'd81,  12'd399,  12'd204,  -12'd50,  12'd255,  -12'd13,  12'd226,  -12'd194,  12'd278,  -12'd95,  12'd370,  -12'd355,  -12'd150,  -12'd340,  12'd97,  -12'd8,  
12'd26,  -12'd62,  -12'd308,  12'd364,  -12'd73,  12'd46,  12'd52,  -12'd401,  -12'd102,  12'd369,  -12'd133,  -12'd136,  -12'd46,  -12'd318,  12'd169,  12'd30,  
-12'd416,  -12'd70,  12'd319,  12'd244,  12'd81,  -12'd229,  -12'd18,  12'd119,  -12'd183,  12'd182,  -12'd86,  12'd390,  -12'd158,  12'd243,  -12'd320,  12'd31,  
12'd180,  -12'd37,  -12'd312,  -12'd40,  -12'd185,  -12'd146,  -12'd442,  -12'd265,  -12'd311,  12'd321,  -12'd67,  12'd13,  12'd20,  12'd645,  -12'd261,  -12'd99,  
12'd7,  12'd209,  -12'd210,  12'd64,  -12'd108,  -12'd97,  -12'd498,  -12'd6,  12'd116,  -12'd160,  -12'd272,  -12'd187,  12'd14,  12'd92,  12'd86,  -12'd143,  
12'd238,  -12'd38,  -12'd503,  -12'd132,  -12'd138,  12'd228,  -12'd12,  12'd264,  -12'd138,  -12'd451,  12'd260,  -12'd125,  -12'd151,  -12'd176,  12'd186,  12'd158,  
12'd267,  12'd169,  -12'd127,  12'd158,  -12'd154,  12'd30,  -12'd145,  12'd193,  12'd16,  -12'd398,  12'd35,  12'd107,  12'd108,  -12'd13,  -12'd56,  12'd63,  
-12'd320,  -12'd157,  -12'd396,  -12'd117,  -12'd108,  -12'd135,  12'd62,  12'd67,  -12'd391,  -12'd835,  -12'd167,  -12'd426,  -12'd325,  -12'd39,  -12'd38,  -12'd223,  

12'd222,  12'd202,  12'd449,  12'd314,  12'd212,  12'd78,  12'd275,  12'd137,  12'd315,  12'd227,  12'd144,  -12'd173,  12'd161,  12'd479,  12'd272,  -12'd387,  
-12'd363,  -12'd370,  12'd266,  12'd269,  12'd244,  -12'd1,  -12'd155,  -12'd167,  -12'd127,  12'd298,  12'd62,  12'd81,  -12'd31,  -12'd40,  -12'd32,  12'd43,  
-12'd153,  -12'd16,  -12'd26,  12'd74,  -12'd175,  12'd156,  12'd69,  12'd148,  12'd12,  12'd47,  12'd273,  12'd401,  12'd51,  -12'd630,  -12'd120,  -12'd416,  
12'd199,  -12'd24,  -12'd36,  -12'd72,  12'd408,  -12'd313,  -12'd327,  12'd38,  -12'd221,  12'd285,  -12'd16,  -12'd230,  12'd311,  -12'd676,  -12'd421,  12'd294,  
12'd383,  -12'd436,  -12'd384,  -12'd12,  -12'd248,  12'd29,  -12'd273,  12'd376,  -12'd87,  12'd90,  -12'd128,  -12'd412,  -12'd63,  -12'd233,  -12'd91,  -12'd119,  
-12'd177,  12'd282,  -12'd291,  12'd284,  12'd228,  12'd101,  -12'd253,  12'd313,  12'd141,  12'd149,  12'd322,  12'd67,  -12'd76,  -12'd25,  12'd436,  -12'd89,  
-12'd93,  -12'd115,  12'd132,  12'd184,  12'd151,  12'd139,  12'd44,  12'd162,  12'd126,  12'd213,  12'd100,  12'd198,  -12'd171,  -12'd287,  -12'd132,  -12'd217,  
-12'd664,  12'd242,  -12'd387,  -12'd145,  12'd312,  -12'd381,  12'd262,  12'd300,  -12'd31,  12'd10,  12'd134,  12'd79,  12'd59,  -12'd77,  12'd97,  -12'd42,  
12'd152,  12'd11,  -12'd5,  12'd181,  12'd92,  -12'd21,  -12'd381,  -12'd46,  -12'd248,  12'd75,  12'd2,  -12'd3,  12'd151,  -12'd3,  12'd104,  -12'd20,  
12'd476,  -12'd112,  -12'd458,  -12'd8,  -12'd185,  12'd3,  -12'd215,  12'd9,  12'd22,  12'd363,  12'd163,  12'd105,  12'd273,  -12'd490,  12'd131,  12'd273,  
12'd161,  12'd42,  -12'd88,  12'd95,  12'd426,  -12'd174,  -12'd111,  12'd42,  -12'd184,  -12'd422,  12'd205,  12'd90,  12'd51,  -12'd9,  -12'd61,  -12'd108,  
-12'd4,  12'd30,  -12'd57,  -12'd242,  -12'd254,  -12'd136,  -12'd229,  -12'd369,  -12'd68,  -12'd7,  12'd402,  -12'd51,  12'd18,  -12'd385,  12'd268,  12'd99,  
12'd34,  -12'd182,  12'd138,  12'd120,  -12'd246,  -12'd122,  -12'd116,  12'd155,  -12'd38,  -12'd259,  12'd684,  -12'd257,  -12'd126,  12'd327,  12'd358,  12'd122,  
-12'd31,  12'd210,  12'd53,  12'd273,  12'd57,  12'd13,  12'd67,  -12'd1,  12'd288,  -12'd324,  12'd66,  12'd106,  12'd311,  -12'd113,  -12'd71,  12'd191,  
-12'd613,  -12'd225,  12'd178,  12'd447,  12'd126,  12'd168,  12'd6,  -12'd107,  12'd104,  12'd130,  12'd219,  12'd65,  12'd381,  12'd57,  12'd354,  -12'd83,  
12'd193,  12'd134,  12'd78,  -12'd141,  12'd104,  -12'd239,  12'd60,  12'd115,  -12'd270,  -12'd28,  12'd306,  12'd14,  12'd190,  -12'd129,  12'd14,  -12'd66,  
-12'd198,  12'd35,  -12'd426,  -12'd314,  -12'd52,  -12'd485,  -12'd41,  -12'd146,  -12'd82,  -12'd76,  12'd133,  12'd61,  12'd67,  12'd51,  -12'd454,  12'd180,  
12'd289,  12'd374,  12'd3,  -12'd411,  12'd66,  -12'd339,  12'd83,  -12'd25,  12'd97,  12'd208,  -12'd11,  -12'd144,  -12'd103,  12'd319,  -12'd31,  -12'd22,  
12'd345,  12'd453,  12'd411,  -12'd289,  -12'd2,  -12'd66,  12'd71,  12'd300,  12'd376,  12'd138,  12'd160,  12'd302,  -12'd310,  -12'd26,  12'd368,  -12'd205,  
12'd69,  12'd177,  -12'd28,  12'd263,  12'd344,  12'd114,  -12'd43,  12'd58,  12'd129,  -12'd30,  12'd335,  -12'd363,  12'd34,  12'd183,  -12'd134,  12'd310,  
-12'd10,  12'd42,  -12'd105,  -12'd440,  12'd12,  -12'd136,  12'd216,  -12'd409,  12'd81,  -12'd521,  -12'd343,  12'd146,  -12'd515,  -12'd396,  12'd51,  12'd170,  
-12'd140,  -12'd85,  -12'd450,  -12'd33,  -12'd13,  -12'd51,  12'd318,  -12'd197,  12'd399,  -12'd192,  -12'd253,  12'd131,  -12'd175,  12'd75,  -12'd102,  12'd15,  
12'd254,  -12'd158,  12'd305,  -12'd121,  12'd189,  -12'd52,  12'd338,  -12'd317,  12'd774,  12'd91,  -12'd48,  -12'd26,  -12'd223,  12'd263,  -12'd115,  -12'd280,  
-12'd148,  12'd86,  12'd158,  -12'd177,  -12'd5,  -12'd161,  -12'd203,  12'd215,  12'd6,  12'd8,  -12'd236,  -12'd196,  -12'd16,  12'd334,  12'd37,  -12'd138,  
-12'd210,  12'd59,  12'd106,  12'd116,  -12'd238,  12'd58,  -12'd210,  -12'd20,  12'd99,  12'd473,  12'd66,  -12'd83,  -12'd307,  -12'd105,  -12'd366,  -12'd87,  

12'd99,  12'd459,  12'd125,  -12'd104,  -12'd181,  12'd26,  12'd580,  -12'd141,  12'd26,  -12'd29,  -12'd34,  12'd532,  -12'd430,  12'd398,  -12'd407,  12'd81,  
12'd5,  12'd190,  -12'd199,  -12'd112,  -12'd414,  -12'd156,  12'd497,  12'd56,  12'd274,  -12'd82,  -12'd49,  12'd42,  -12'd307,  12'd1,  12'd88,  12'd68,  
12'd430,  12'd152,  -12'd7,  -12'd289,  12'd209,  -12'd249,  -12'd97,  12'd153,  12'd265,  -12'd3,  12'd19,  12'd13,  12'd97,  12'd23,  12'd11,  -12'd130,  
-12'd18,  -12'd57,  12'd22,  12'd84,  -12'd27,  12'd339,  12'd130,  12'd11,  12'd133,  12'd134,  -12'd100,  -12'd171,  12'd244,  -12'd184,  -12'd64,  -12'd1,  
-12'd538,  12'd376,  12'd197,  -12'd70,  -12'd269,  12'd269,  -12'd129,  12'd13,  12'd109,  -12'd77,  12'd362,  12'd18,  12'd265,  12'd388,  12'd309,  12'd342,  
-12'd290,  -12'd359,  12'd65,  -12'd276,  -12'd200,  -12'd104,  12'd290,  12'd80,  12'd255,  -12'd121,  -12'd35,  -12'd98,  -12'd351,  12'd93,  12'd129,  12'd76,  
12'd223,  -12'd84,  12'd107,  -12'd387,  12'd101,  12'd32,  -12'd291,  -12'd154,  12'd229,  12'd111,  -12'd159,  -12'd113,  -12'd93,  12'd295,  12'd198,  12'd16,  
-12'd287,  -12'd219,  -12'd9,  -12'd215,  12'd114,  -12'd133,  12'd60,  12'd263,  -12'd156,  12'd176,  12'd269,  12'd145,  -12'd426,  -12'd138,  12'd43,  -12'd200,  
-12'd70,  -12'd14,  -12'd17,  -12'd134,  12'd224,  12'd47,  -12'd75,  -12'd159,  -12'd219,  12'd568,  -12'd95,  -12'd14,  12'd22,  -12'd252,  12'd33,  -12'd59,  
-12'd321,  -12'd287,  -12'd81,  -12'd81,  -12'd270,  -12'd362,  12'd203,  12'd71,  12'd29,  12'd125,  -12'd151,  -12'd106,  -12'd160,  -12'd139,  -12'd428,  12'd207,  
-12'd164,  12'd245,  -12'd73,  -12'd22,  12'd78,  12'd341,  -12'd180,  12'd74,  -12'd379,  12'd410,  -12'd261,  -12'd69,  12'd35,  -12'd17,  12'd99,  12'd54,  
12'd473,  12'd188,  12'd71,  12'd39,  -12'd23,  12'd107,  -12'd1,  12'd245,  -12'd34,  -12'd81,  12'd133,  -12'd212,  -12'd474,  12'd417,  12'd64,  -12'd360,  
-12'd106,  12'd236,  -12'd215,  -12'd19,  12'd386,  12'd143,  12'd85,  12'd150,  12'd376,  -12'd180,  -12'd98,  12'd341,  -12'd199,  -12'd227,  -12'd169,  -12'd288,  
12'd72,  12'd68,  -12'd279,  -12'd608,  12'd224,  12'd194,  12'd115,  -12'd279,  12'd414,  12'd271,  -12'd101,  -12'd268,  12'd30,  -12'd27,  -12'd64,  -12'd73,  
-12'd332,  -12'd205,  -12'd196,  12'd297,  -12'd417,  12'd263,  -12'd255,  -12'd78,  12'd200,  12'd271,  12'd97,  -12'd26,  -12'd435,  -12'd39,  -12'd37,  12'd385,  
12'd52,  -12'd48,  12'd374,  12'd191,  -12'd39,  12'd77,  -12'd34,  -12'd68,  -12'd183,  -12'd78,  -12'd442,  12'd277,  -12'd144,  12'd122,  -12'd6,  12'd181,  
12'd296,  12'd89,  -12'd191,  12'd327,  -12'd67,  12'd104,  -12'd199,  12'd54,  12'd471,  -12'd176,  -12'd301,  12'd175,  12'd221,  12'd152,  12'd393,  12'd144,  
-12'd166,  -12'd158,  -12'd19,  12'd31,  -12'd45,  12'd88,  12'd331,  12'd390,  -12'd288,  -12'd296,  12'd4,  -12'd77,  -12'd473,  12'd194,  12'd231,  -12'd63,  
-12'd19,  12'd152,  -12'd136,  12'd39,  12'd211,  12'd155,  -12'd74,  -12'd363,  -12'd135,  -12'd53,  -12'd213,  12'd273,  -12'd14,  12'd499,  12'd21,  -12'd187,  
-12'd179,  12'd134,  12'd322,  12'd126,  -12'd102,  12'd160,  12'd291,  -12'd238,  12'd321,  12'd48,  -12'd103,  -12'd11,  -12'd257,  12'd242,  -12'd103,  -12'd38,  
-12'd406,  -12'd281,  -12'd152,  12'd246,  12'd185,  12'd504,  -12'd181,  12'd487,  12'd149,  12'd73,  -12'd197,  -12'd218,  12'd255,  -12'd288,  12'd16,  12'd163,  
12'd14,  12'd293,  12'd43,  12'd186,  12'd567,  -12'd3,  -12'd253,  12'd516,  -12'd166,  -12'd273,  12'd448,  -12'd225,  -12'd6,  -12'd205,  12'd339,  -12'd9,  
-12'd172,  -12'd175,  -12'd209,  12'd305,  12'd31,  12'd309,  -12'd98,  12'd334,  12'd111,  12'd280,  12'd267,  12'd48,  12'd249,  -12'd52,  12'd18,  12'd126,  
12'd21,  12'd356,  -12'd273,  12'd415,  -12'd104,  12'd397,  12'd1,  12'd176,  12'd64,  12'd285,  -12'd265,  12'd524,  12'd338,  -12'd30,  12'd32,  -12'd130,  
12'd488,  12'd110,  12'd163,  12'd379,  12'd149,  12'd72,  12'd128,  12'd431,  12'd695,  12'd108,  12'd180,  12'd349,  -12'd12,  12'd243,  -12'd77,  -12'd80,  

-12'd79,  -12'd42,  12'd86,  12'd36,  -12'd41,  12'd116,  12'd353,  12'd246,  -12'd314,  -12'd191,  -12'd61,  -12'd30,  -12'd93,  -12'd288,  12'd41,  -12'd80,  
12'd49,  -12'd319,  12'd33,  -12'd276,  12'd86,  -12'd54,  -12'd258,  -12'd432,  -12'd407,  -12'd210,  -12'd126,  -12'd280,  12'd37,  12'd60,  -12'd401,  -12'd307,  
-12'd16,  12'd59,  12'd116,  12'd187,  -12'd298,  -12'd104,  -12'd181,  -12'd58,  -12'd19,  12'd44,  -12'd32,  -12'd480,  12'd20,  12'd168,  -12'd272,  12'd210,  
-12'd319,  -12'd152,  -12'd311,  12'd68,  12'd122,  -12'd386,  -12'd43,  -12'd147,  12'd74,  -12'd188,  -12'd87,  12'd43,  -12'd46,  12'd14,  -12'd66,  -12'd30,  
-12'd21,  12'd60,  -12'd234,  -12'd202,  12'd4,  -12'd73,  -12'd73,  12'd33,  12'd66,  12'd243,  -12'd171,  12'd32,  12'd61,  -12'd165,  -12'd258,  -12'd258,  
-12'd162,  -12'd147,  -12'd93,  -12'd162,  -12'd384,  12'd262,  -12'd249,  12'd225,  12'd228,  -12'd10,  -12'd182,  -12'd273,  12'd248,  -12'd118,  12'd199,  -12'd290,  
-12'd16,  12'd26,  12'd10,  12'd223,  12'd168,  12'd260,  -12'd271,  -12'd453,  -12'd68,  12'd273,  12'd241,  -12'd113,  12'd150,  12'd150,  12'd151,  -12'd303,  
12'd280,  12'd175,  -12'd166,  -12'd342,  12'd95,  12'd150,  -12'd47,  12'd62,  -12'd109,  -12'd20,  -12'd261,  12'd101,  12'd104,  12'd147,  -12'd198,  -12'd265,  
-12'd135,  -12'd47,  -12'd257,  12'd0,  12'd32,  -12'd226,  -12'd298,  -12'd269,  -12'd99,  12'd71,  -12'd246,  -12'd85,  -12'd272,  -12'd81,  12'd92,  -12'd126,  
12'd272,  12'd113,  12'd343,  -12'd209,  -12'd184,  12'd161,  -12'd114,  -12'd110,  -12'd202,  12'd138,  -12'd117,  -12'd330,  -12'd304,  12'd150,  -12'd253,  12'd85,  
-12'd188,  -12'd267,  -12'd294,  12'd59,  -12'd158,  12'd107,  -12'd154,  -12'd407,  12'd194,  -12'd198,  -12'd411,  -12'd66,  -12'd84,  -12'd70,  -12'd70,  -12'd210,  
12'd88,  -12'd193,  -12'd15,  -12'd97,  -12'd326,  -12'd74,  12'd91,  -12'd187,  -12'd190,  12'd169,  -12'd147,  -12'd243,  -12'd249,  -12'd154,  12'd121,  -12'd210,  
12'd107,  -12'd55,  -12'd354,  12'd113,  -12'd138,  -12'd396,  -12'd9,  12'd127,  -12'd76,  -12'd182,  12'd61,  -12'd425,  -12'd159,  -12'd97,  12'd206,  -12'd14,  
12'd88,  -12'd272,  -12'd365,  12'd305,  -12'd174,  -12'd35,  -12'd38,  -12'd159,  -12'd394,  12'd4,  -12'd226,  -12'd308,  -12'd132,  -12'd61,  12'd222,  -12'd60,  
12'd126,  12'd83,  -12'd240,  12'd84,  -12'd5,  -12'd90,  -12'd192,  -12'd33,  -12'd230,  12'd207,  -12'd112,  -12'd95,  12'd53,  12'd344,  -12'd137,  12'd255,  
-12'd3,  12'd104,  -12'd221,  -12'd173,  -12'd64,  -12'd85,  12'd63,  -12'd98,  12'd116,  -12'd249,  12'd186,  -12'd130,  -12'd210,  12'd1,  -12'd113,  -12'd48,  
12'd216,  -12'd227,  12'd122,  -12'd8,  -12'd312,  -12'd276,  -12'd66,  12'd38,  -12'd12,  -12'd396,  -12'd134,  12'd101,  -12'd7,  -12'd120,  -12'd463,  -12'd144,  
12'd232,  -12'd127,  -12'd282,  -12'd205,  12'd144,  -12'd179,  -12'd145,  -12'd135,  12'd65,  -12'd411,  -12'd215,  -12'd70,  12'd130,  -12'd430,  12'd169,  12'd83,  
12'd10,  -12'd147,  12'd84,  -12'd95,  -12'd26,  12'd243,  12'd144,  -12'd233,  -12'd195,  12'd90,  -12'd124,  12'd16,  12'd40,  -12'd121,  -12'd346,  -12'd194,  
12'd26,  -12'd101,  -12'd205,  -12'd418,  12'd117,  12'd122,  -12'd417,  -12'd437,  -12'd21,  12'd178,  -12'd41,  12'd173,  -12'd340,  -12'd11,  12'd5,  12'd49,  
-12'd140,  -12'd228,  -12'd449,  -12'd115,  -12'd360,  -12'd388,  -12'd75,  -12'd373,  -12'd290,  -12'd212,  -12'd43,  -12'd84,  -12'd146,  12'd200,  -12'd159,  -12'd52,  
-12'd241,  12'd37,  -12'd71,  -12'd409,  -12'd292,  -12'd291,  12'd53,  -12'd309,  12'd144,  -12'd147,  -12'd236,  12'd63,  -12'd218,  -12'd133,  -12'd417,  12'd7,  
12'd254,  -12'd85,  -12'd58,  12'd93,  -12'd18,  -12'd42,  -12'd179,  12'd41,  12'd172,  12'd9,  -12'd111,  -12'd357,  -12'd28,  -12'd264,  12'd15,  -12'd18,  
12'd326,  12'd126,  12'd202,  -12'd385,  -12'd84,  12'd36,  -12'd267,  -12'd139,  -12'd304,  12'd164,  -12'd385,  12'd52,  -12'd374,  12'd157,  -12'd319,  -12'd123,  
12'd341,  12'd262,  -12'd42,  -12'd239,  -12'd90,  -12'd252,  12'd82,  -12'd11,  12'd117,  -12'd11,  12'd305,  -12'd273,  -12'd85,  12'd22,  -12'd7,  -12'd261,  

12'd147,  -12'd342,  12'd184,  -12'd149,  -12'd263,  -12'd51,  -12'd209,  -12'd164,  -12'd31,  12'd441,  -12'd369,  -12'd379,  -12'd385,  -12'd161,  -12'd488,  -12'd100,  
-12'd260,  -12'd571,  -12'd154,  -12'd12,  -12'd68,  12'd307,  12'd32,  -12'd1,  -12'd555,  -12'd0,  -12'd312,  -12'd461,  -12'd296,  -12'd557,  -12'd270,  12'd56,  
-12'd109,  12'd150,  -12'd12,  12'd167,  -12'd346,  12'd123,  -12'd591,  -12'd132,  -12'd102,  -12'd228,  -12'd518,  12'd140,  -12'd120,  12'd67,  -12'd442,  -12'd197,  
-12'd69,  12'd195,  -12'd10,  12'd30,  12'd57,  12'd473,  -12'd123,  -12'd311,  12'd166,  -12'd106,  -12'd309,  -12'd295,  -12'd249,  -12'd374,  -12'd81,  12'd109,  
12'd443,  12'd323,  12'd175,  12'd336,  -12'd273,  12'd191,  -12'd127,  12'd188,  12'd215,  -12'd163,  -12'd64,  -12'd327,  -12'd154,  -12'd138,  12'd56,  12'd116,  
-12'd369,  -12'd240,  -12'd526,  12'd52,  -12'd142,  -12'd258,  -12'd546,  -12'd365,  -12'd104,  12'd177,  12'd458,  12'd372,  12'd52,  -12'd68,  -12'd67,  -12'd301,  
-12'd137,  -12'd178,  12'd48,  12'd211,  12'd44,  12'd186,  -12'd153,  -12'd253,  12'd218,  12'd186,  12'd481,  -12'd266,  12'd184,  -12'd47,  -12'd28,  -12'd0,  
12'd253,  12'd107,  12'd99,  12'd261,  12'd37,  12'd132,  -12'd27,  12'd442,  12'd58,  12'd217,  -12'd2,  -12'd40,  12'd408,  12'd345,  12'd84,  -12'd53,  
12'd508,  12'd5,  -12'd46,  -12'd67,  12'd134,  12'd355,  -12'd165,  12'd70,  12'd401,  -12'd52,  12'd635,  -12'd149,  12'd185,  12'd246,  -12'd63,  -12'd1,  
12'd114,  12'd134,  12'd149,  -12'd68,  12'd410,  -12'd341,  -12'd353,  -12'd27,  -12'd134,  12'd542,  -12'd393,  12'd256,  -12'd153,  12'd463,  12'd0,  12'd120,  
-12'd340,  12'd55,  -12'd439,  12'd39,  -12'd123,  12'd221,  12'd361,  12'd126,  12'd599,  -12'd94,  12'd421,  -12'd298,  -12'd20,  12'd175,  12'd356,  12'd304,  
-12'd168,  12'd21,  -12'd136,  12'd85,  -12'd27,  -12'd150,  12'd102,  -12'd307,  12'd360,  -12'd25,  12'd243,  -12'd237,  -12'd460,  12'd481,  12'd414,  12'd273,  
-12'd105,  -12'd188,  -12'd175,  -12'd259,  12'd28,  -12'd477,  -12'd214,  12'd137,  -12'd458,  -12'd105,  -12'd161,  -12'd462,  -12'd55,  12'd115,  12'd371,  12'd286,  
12'd108,  12'd162,  -12'd265,  -12'd107,  -12'd192,  -12'd294,  -12'd526,  -12'd81,  -12'd259,  -12'd93,  12'd10,  -12'd210,  -12'd482,  12'd334,  12'd89,  12'd69,  
12'd261,  -12'd83,  12'd401,  -12'd176,  -12'd197,  -12'd288,  12'd37,  -12'd406,  12'd147,  12'd465,  -12'd409,  12'd412,  -12'd319,  12'd99,  12'd97,  12'd168,  
-12'd67,  -12'd467,  12'd309,  -12'd37,  -12'd152,  -12'd189,  12'd50,  -12'd116,  -12'd322,  12'd39,  12'd446,  -12'd344,  -12'd354,  -12'd352,  -12'd340,  -12'd29,  
12'd121,  -12'd180,  -12'd217,  12'd156,  -12'd253,  -12'd352,  -12'd142,  12'd52,  -12'd421,  -12'd386,  12'd89,  -12'd419,  -12'd20,  -12'd78,  -12'd258,  12'd63,  
12'd47,  12'd388,  -12'd115,  -12'd27,  -12'd285,  -12'd164,  12'd199,  12'd138,  12'd505,  12'd250,  -12'd270,  -12'd238,  -12'd422,  -12'd155,  -12'd192,  -12'd306,  
12'd114,  12'd238,  12'd51,  -12'd210,  -12'd440,  12'd69,  12'd24,  12'd146,  12'd146,  12'd13,  12'd30,  12'd176,  -12'd223,  12'd127,  -12'd72,  -12'd245,  
12'd389,  -12'd117,  12'd119,  -12'd60,  -12'd333,  12'd301,  12'd110,  12'd255,  12'd201,  -12'd45,  12'd226,  12'd40,  12'd313,  12'd212,  12'd322,  12'd116,  
-12'd390,  12'd428,  -12'd496,  -12'd382,  12'd282,  -12'd304,  -12'd458,  -12'd391,  -12'd153,  -12'd371,  -12'd230,  12'd163,  -12'd81,  12'd182,  -12'd160,  -12'd76,  
-12'd85,  12'd171,  12'd85,  -12'd606,  -12'd79,  -12'd277,  -12'd214,  -12'd373,  -12'd355,  -12'd165,  12'd87,  -12'd55,  -12'd292,  12'd79,  -12'd7,  -12'd324,  
12'd292,  -12'd199,  12'd340,  -12'd28,  -12'd289,  -12'd182,  -12'd241,  -12'd53,  12'd343,  -12'd57,  -12'd568,  -12'd7,  -12'd474,  12'd31,  12'd139,  -12'd337,  
12'd471,  -12'd443,  12'd260,  12'd6,  12'd265,  12'd78,  -12'd150,  -12'd255,  12'd19,  12'd355,  12'd146,  -12'd6,  12'd79,  12'd57,  12'd74,  -12'd9,  
12'd292,  -12'd170,  -12'd371,  -12'd69,  12'd68,  12'd280,  -12'd15,  12'd258,  12'd171,  -12'd1,  12'd155,  12'd157,  -12'd17,  -12'd175,  12'd530,  12'd269,  

-12'd66,  -12'd293,  -12'd131,  12'd461,  12'd91,  12'd333,  12'd154,  12'd294,  12'd233,  12'd172,  12'd408,  -12'd7,  12'd213,  -12'd144,  12'd147,  -12'd4,  
-12'd403,  -12'd202,  12'd345,  12'd427,  12'd40,  12'd208,  -12'd164,  12'd272,  12'd104,  12'd480,  12'd349,  -12'd307,  12'd286,  -12'd120,  12'd489,  -12'd186,  
-12'd207,  -12'd454,  -12'd102,  -12'd1,  -12'd317,  12'd62,  -12'd218,  12'd242,  -12'd31,  12'd60,  -12'd54,  12'd85,  12'd347,  -12'd746,  -12'd108,  -12'd76,  
12'd192,  12'd91,  -12'd44,  12'd169,  12'd151,  12'd138,  -12'd189,  -12'd137,  -12'd158,  12'd26,  -12'd227,  12'd189,  12'd377,  -12'd755,  -12'd151,  -12'd51,  
-12'd17,  12'd78,  12'd45,  12'd65,  -12'd138,  12'd102,  -12'd127,  -12'd61,  -12'd235,  -12'd233,  -12'd290,  -12'd82,  12'd469,  -12'd76,  -12'd27,  12'd145,  
-12'd163,  -12'd213,  -12'd165,  12'd137,  -12'd97,  -12'd140,  -12'd516,  12'd64,  -12'd104,  -12'd131,  12'd247,  12'd3,  12'd30,  12'd346,  12'd90,  -12'd48,  
-12'd74,  12'd85,  -12'd93,  12'd123,  12'd6,  12'd49,  -12'd42,  -12'd53,  12'd224,  -12'd336,  12'd90,  12'd125,  12'd170,  12'd188,  -12'd57,  -12'd133,  
-12'd485,  12'd221,  -12'd97,  12'd88,  -12'd233,  12'd172,  -12'd390,  -12'd142,  12'd704,  12'd45,  12'd178,  12'd42,  12'd37,  -12'd307,  -12'd76,  12'd178,  
-12'd31,  -12'd133,  -12'd344,  -12'd71,  -12'd236,  -12'd209,  -12'd415,  12'd211,  12'd212,  12'd404,  -12'd139,  12'd144,  12'd436,  -12'd581,  -12'd153,  12'd259,  
12'd129,  12'd50,  -12'd250,  -12'd50,  12'd391,  12'd65,  12'd126,  12'd128,  12'd222,  12'd150,  12'd273,  -12'd149,  12'd50,  -12'd97,  -12'd372,  12'd132,  
-12'd118,  -12'd10,  12'd303,  12'd87,  -12'd171,  12'd150,  -12'd41,  12'd204,  12'd0,  -12'd44,  -12'd79,  -12'd323,  12'd103,  12'd104,  -12'd341,  12'd97,  
12'd89,  12'd3,  12'd381,  -12'd129,  -12'd80,  -12'd197,  12'd286,  12'd120,  -12'd170,  -12'd342,  12'd235,  -12'd210,  -12'd148,  -12'd160,  12'd196,  12'd118,  
12'd162,  12'd78,  12'd141,  -12'd186,  -12'd257,  -12'd93,  12'd138,  -12'd91,  -12'd184,  12'd50,  -12'd38,  -12'd313,  -12'd9,  12'd18,  -12'd58,  12'd435,  
-12'd264,  12'd312,  -12'd46,  12'd65,  12'd44,  12'd322,  -12'd38,  12'd206,  12'd261,  12'd18,  -12'd88,  -12'd119,  12'd120,  -12'd33,  12'd124,  12'd250,  
-12'd787,  -12'd98,  -12'd255,  -12'd83,  -12'd28,  -12'd449,  12'd90,  12'd25,  12'd59,  -12'd56,  12'd414,  12'd197,  -12'd266,  -12'd111,  12'd386,  12'd116,  
12'd69,  -12'd34,  12'd7,  -12'd74,  -12'd288,  -12'd156,  12'd285,  -12'd426,  12'd226,  -12'd11,  12'd107,  -12'd98,  -12'd56,  12'd46,  -12'd367,  -12'd385,  
-12'd157,  -12'd140,  -12'd180,  -12'd243,  -12'd117,  12'd66,  -12'd141,  12'd209,  -12'd339,  12'd510,  12'd356,  12'd162,  -12'd127,  12'd0,  -12'd1,  12'd46,  
-12'd26,  12'd94,  -12'd181,  12'd169,  12'd70,  12'd2,  -12'd300,  12'd232,  12'd219,  -12'd250,  -12'd200,  -12'd106,  12'd66,  12'd276,  -12'd4,  -12'd362,  
12'd75,  -12'd41,  12'd307,  -12'd52,  12'd107,  12'd92,  -12'd0,  -12'd89,  -12'd254,  -12'd205,  12'd232,  12'd12,  -12'd274,  -12'd56,  -12'd265,  -12'd191,  
12'd163,  12'd300,  12'd241,  -12'd181,  -12'd20,  -12'd70,  12'd188,  12'd272,  12'd47,  -12'd8,  12'd120,  -12'd10,  -12'd109,  12'd304,  -12'd56,  -12'd336,  
12'd147,  -12'd80,  -12'd51,  12'd324,  -12'd283,  -12'd313,  12'd460,  12'd15,  12'd481,  12'd135,  12'd132,  12'd47,  -12'd162,  -12'd501,  12'd14,  12'd263,  
-12'd124,  12'd7,  -12'd363,  12'd281,  -12'd105,  12'd82,  12'd222,  -12'd72,  12'd105,  -12'd166,  12'd7,  -12'd74,  -12'd160,  12'd115,  -12'd302,  12'd230,  
12'd176,  -12'd81,  12'd289,  -12'd292,  -12'd42,  -12'd196,  -12'd53,  12'd112,  12'd556,  -12'd52,  12'd175,  12'd45,  -12'd81,  12'd54,  -12'd370,  -12'd218,  
12'd117,  12'd340,  12'd57,  12'd142,  -12'd165,  -12'd87,  -12'd23,  -12'd36,  12'd444,  -12'd35,  12'd156,  -12'd271,  12'd129,  12'd101,  -12'd23,  -12'd51,  
12'd71,  12'd158,  -12'd50,  -12'd461,  -12'd298,  -12'd262,  -12'd65,  -12'd30,  -12'd15,  -12'd237,  -12'd233,  -12'd250,  -12'd106,  12'd207,  -12'd102,  -12'd120,  

-12'd346,  12'd119,  12'd300,  12'd405,  12'd26,  12'd131,  -12'd596,  12'd592,  -12'd123,  12'd553,  -12'd499,  12'd60,  12'd242,  -12'd205,  -12'd60,  -12'd20,  
-12'd14,  12'd238,  12'd872,  12'd139,  12'd328,  -12'd33,  -12'd45,  12'd270,  12'd280,  -12'd12,  -12'd210,  -12'd96,  -12'd88,  12'd483,  -12'd138,  -12'd386,  
12'd173,  12'd72,  12'd741,  12'd173,  -12'd350,  12'd100,  12'd261,  -12'd153,  12'd58,  -12'd246,  -12'd51,  -12'd72,  -12'd152,  12'd510,  12'd200,  -12'd327,  
12'd52,  -12'd2,  12'd71,  12'd307,  -12'd79,  -12'd257,  12'd127,  12'd119,  -12'd207,  -12'd4,  12'd360,  12'd220,  12'd280,  -12'd174,  -12'd244,  -12'd258,  
12'd271,  12'd536,  -12'd215,  -12'd26,  -12'd168,  12'd391,  12'd129,  -12'd94,  12'd245,  12'd123,  12'd269,  -12'd190,  12'd299,  12'd218,  -12'd93,  12'd167,  
-12'd93,  12'd420,  12'd447,  12'd14,  12'd333,  12'd406,  -12'd387,  12'd63,  -12'd140,  12'd44,  -12'd267,  -12'd67,  12'd259,  12'd172,  12'd75,  12'd208,  
12'd296,  12'd76,  12'd348,  12'd298,  -12'd69,  12'd241,  -12'd189,  -12'd40,  12'd407,  -12'd43,  -12'd156,  12'd138,  -12'd86,  12'd203,  12'd27,  -12'd34,  
12'd199,  12'd177,  12'd591,  12'd344,  -12'd133,  12'd1,  -12'd300,  12'd63,  -12'd98,  -12'd5,  12'd249,  -12'd156,  -12'd382,  12'd371,  12'd141,  -12'd117,  
12'd9,  12'd286,  12'd502,  -12'd326,  -12'd174,  12'd25,  12'd33,  -12'd86,  -12'd67,  -12'd181,  -12'd206,  12'd50,  12'd93,  12'd189,  -12'd188,  -12'd135,  
12'd126,  12'd62,  -12'd265,  12'd281,  12'd4,  -12'd405,  -12'd67,  -12'd95,  12'd155,  -12'd152,  12'd412,  -12'd171,  -12'd84,  12'd56,  -12'd236,  12'd7,  
-12'd301,  12'd82,  -12'd269,  12'd248,  12'd195,  12'd88,  -12'd124,  12'd300,  12'd213,  12'd140,  12'd380,  12'd161,  12'd220,  12'd7,  12'd123,  12'd145,  
-12'd49,  -12'd200,  -12'd1,  12'd172,  12'd331,  -12'd33,  12'd329,  -12'd75,  12'd309,  12'd36,  -12'd248,  -12'd208,  12'd86,  -12'd29,  12'd249,  12'd269,  
-12'd199,  12'd161,  12'd487,  -12'd182,  -12'd68,  12'd43,  -12'd179,  12'd221,  -12'd80,  -12'd233,  -12'd48,  12'd81,  -12'd28,  12'd240,  -12'd139,  -12'd159,  
-12'd400,  -12'd194,  -12'd430,  12'd251,  -12'd49,  -12'd114,  -12'd100,  12'd219,  -12'd140,  12'd157,  12'd241,  -12'd3,  -12'd317,  -12'd200,  12'd223,  12'd13,  
-12'd450,  12'd40,  12'd362,  12'd153,  -12'd14,  -12'd311,  -12'd26,  12'd57,  -12'd242,  12'd99,  12'd278,  -12'd494,  -12'd147,  -12'd384,  12'd338,  -12'd142,  
-12'd354,  12'd102,  -12'd117,  -12'd84,  -12'd83,  -12'd35,  -12'd120,  -12'd346,  12'd114,  12'd109,  12'd422,  -12'd83,  -12'd9,  -12'd282,  -12'd185,  -12'd37,  
12'd48,  -12'd60,  12'd20,  -12'd0,  12'd176,  12'd89,  -12'd162,  -12'd19,  -12'd63,  12'd514,  -12'd276,  -12'd123,  -12'd115,  12'd205,  -12'd239,  -12'd42,  
-12'd475,  12'd31,  12'd87,  -12'd73,  12'd104,  -12'd225,  -12'd272,  12'd80,  -12'd245,  12'd108,  -12'd451,  -12'd70,  12'd180,  12'd352,  12'd273,  -12'd221,  
-12'd276,  12'd57,  12'd3,  -12'd92,  -12'd409,  -12'd58,  12'd279,  -12'd247,  -12'd95,  -12'd152,  12'd131,  12'd199,  -12'd346,  -12'd353,  -12'd78,  -12'd8,  
12'd188,  12'd200,  12'd523,  -12'd399,  12'd43,  12'd300,  -12'd105,  12'd147,  -12'd100,  12'd106,  12'd240,  12'd481,  -12'd42,  12'd76,  -12'd267,  -12'd49,  
-12'd228,  -12'd120,  -12'd174,  -12'd307,  -12'd108,  12'd73,  12'd53,  -12'd28,  -12'd64,  12'd190,  -12'd224,  -12'd303,  -12'd247,  -12'd130,  -12'd83,  12'd141,  
-12'd74,  -12'd241,  12'd74,  12'd25,  -12'd86,  -12'd72,  -12'd168,  -12'd11,  -12'd223,  12'd39,  12'd75,  -12'd297,  -12'd39,  12'd690,  12'd342,  12'd181,  
-12'd167,  12'd71,  12'd368,  -12'd34,  -12'd265,  12'd238,  -12'd168,  -12'd225,  -12'd231,  -12'd240,  -12'd312,  -12'd32,  -12'd135,  -12'd25,  12'd119,  -12'd126,  
12'd281,  12'd272,  12'd91,  -12'd203,  12'd216,  -12'd285,  -12'd18,  -12'd155,  -12'd200,  -12'd351,  12'd505,  -12'd158,  -12'd85,  -12'd27,  -12'd42,  12'd174,  
12'd214,  -12'd92,  -12'd137,  12'd102,  12'd294,  12'd202,  12'd67,  -12'd119,  12'd27,  -12'd471,  -12'd87,  12'd307,  -12'd67,  12'd272,  12'd126,  12'd22,  

12'd127,  12'd409,  12'd219,  -12'd21,  -12'd123,  12'd414,  -12'd643,  12'd217,  12'd323,  12'd114,  12'd108,  -12'd502,  12'd327,  -12'd34,  -12'd20,  12'd316,  
-12'd123,  12'd506,  12'd421,  12'd103,  12'd137,  -12'd57,  -12'd2,  12'd271,  12'd248,  -12'd278,  12'd327,  12'd95,  -12'd110,  12'd9,  12'd457,  -12'd95,  
-12'd12,  12'd70,  12'd71,  -12'd96,  -12'd155,  12'd43,  -12'd48,  -12'd172,  12'd121,  -12'd327,  12'd3,  -12'd1,  -12'd62,  12'd84,  12'd365,  12'd290,  
-12'd139,  -12'd101,  -12'd45,  12'd75,  -12'd422,  12'd567,  12'd133,  12'd237,  -12'd58,  -12'd209,  12'd497,  12'd44,  12'd116,  12'd297,  12'd276,  -12'd151,  
12'd340,  12'd71,  12'd1,  -12'd52,  -12'd422,  12'd267,  12'd29,  -12'd159,  -12'd31,  -12'd370,  -12'd39,  -12'd160,  12'd84,  12'd187,  -12'd340,  12'd21,  
-12'd429,  12'd239,  12'd104,  -12'd546,  12'd471,  -12'd118,  12'd457,  -12'd28,  -12'd24,  12'd253,  -12'd0,  -12'd233,  12'd40,  -12'd105,  -12'd223,  -12'd70,  
-12'd273,  -12'd200,  -12'd91,  -12'd540,  12'd167,  12'd417,  -12'd216,  12'd31,  -12'd122,  -12'd161,  -12'd486,  -12'd264,  12'd80,  12'd167,  -12'd144,  -12'd216,  
12'd112,  -12'd107,  12'd234,  -12'd86,  -12'd433,  -12'd403,  -12'd354,  -12'd327,  -12'd373,  12'd66,  -12'd6,  -12'd13,  -12'd311,  -12'd46,  12'd77,  -12'd201,  
-12'd72,  -12'd31,  -12'd32,  -12'd238,  -12'd464,  12'd172,  -12'd65,  -12'd184,  -12'd15,  -12'd111,  12'd24,  -12'd284,  -12'd408,  12'd105,  -12'd15,  -12'd429,  
-12'd460,  -12'd313,  12'd526,  12'd30,  -12'd299,  -12'd222,  -12'd18,  12'd174,  -12'd315,  12'd93,  12'd38,  -12'd205,  -12'd331,  12'd81,  12'd79,  12'd162,  
-12'd152,  -12'd227,  -12'd215,  -12'd120,  -12'd198,  -12'd177,  12'd121,  12'd144,  12'd390,  -12'd74,  -12'd439,  -12'd260,  -12'd288,  -12'd38,  12'd4,  -12'd102,  
-12'd154,  -12'd323,  12'd22,  12'd320,  -12'd102,  -12'd33,  12'd168,  -12'd273,  -12'd59,  12'd21,  -12'd462,  12'd245,  -12'd21,  -12'd42,  12'd150,  -12'd387,  
12'd27,  -12'd31,  12'd434,  12'd59,  12'd167,  -12'd224,  -12'd247,  -12'd72,  12'd533,  -12'd42,  12'd35,  12'd514,  -12'd59,  12'd502,  -12'd464,  12'd91,  
-12'd388,  -12'd196,  -12'd595,  12'd205,  -12'd28,  12'd84,  12'd108,  -12'd201,  -12'd217,  -12'd331,  12'd349,  12'd164,  12'd66,  12'd257,  -12'd367,  -12'd43,  
12'd206,  -12'd19,  12'd612,  -12'd158,  12'd550,  -12'd175,  -12'd316,  -12'd199,  12'd196,  12'd218,  -12'd60,  12'd327,  12'd296,  12'd17,  -12'd140,  -12'd18,  
12'd412,  12'd190,  12'd114,  -12'd292,  -12'd545,  12'd125,  12'd230,  -12'd265,  12'd39,  12'd176,  -12'd156,  12'd245,  -12'd91,  12'd213,  12'd151,  12'd248,  
12'd289,  -12'd242,  12'd435,  12'd366,  -12'd387,  -12'd247,  12'd142,  12'd169,  12'd26,  -12'd271,  12'd515,  12'd397,  -12'd244,  -12'd172,  12'd115,  12'd138,  
-12'd210,  12'd64,  12'd258,  12'd346,  12'd406,  -12'd227,  12'd202,  -12'd315,  12'd434,  -12'd140,  -12'd108,  12'd150,  12'd70,  -12'd275,  -12'd227,  -12'd138,  
-12'd105,  12'd56,  -12'd624,  12'd22,  12'd75,  -12'd150,  12'd68,  12'd286,  -12'd160,  12'd86,  12'd48,  12'd433,  12'd13,  -12'd115,  12'd109,  12'd146,  
12'd173,  12'd233,  -12'd228,  -12'd433,  -12'd0,  -12'd169,  -12'd39,  -12'd198,  12'd29,  12'd152,  -12'd375,  -12'd124,  12'd227,  12'd309,  12'd432,  12'd228,  
12'd323,  12'd143,  12'd462,  -12'd134,  12'd317,  -12'd30,  -12'd143,  -12'd10,  -12'd283,  12'd38,  -12'd353,  12'd12,  -12'd176,  12'd563,  12'd73,  -12'd187,  
-12'd102,  12'd429,  -12'd7,  -12'd237,  -12'd424,  -12'd27,  12'd36,  -12'd79,  -12'd366,  -12'd20,  12'd300,  -12'd88,  -12'd39,  -12'd540,  12'd363,  -12'd21,  
-12'd399,  12'd141,  -12'd166,  12'd183,  -12'd296,  -12'd107,  -12'd365,  12'd140,  12'd172,  -12'd247,  12'd247,  -12'd162,  12'd88,  12'd1,  12'd130,  -12'd274,  
12'd216,  12'd281,  -12'd1,  -12'd145,  -12'd34,  12'd218,  -12'd157,  -12'd338,  12'd187,  12'd128,  12'd35,  -12'd187,  -12'd93,  12'd37,  12'd269,  -12'd59,  
-12'd207,  12'd183,  -12'd247,  12'd421,  12'd282,  12'd337,  -12'd80,  12'd158,  12'd4,  12'd109,  12'd312,  12'd25,  12'd368,  -12'd125,  12'd73,  12'd73,  

-12'd310,  12'd350,  12'd118,  12'd68,  12'd224,  -12'd45,  -12'd559,  12'd189,  12'd11,  12'd273,  12'd411,  -12'd119,  -12'd57,  -12'd187,  12'd207,  -12'd8,  
-12'd250,  -12'd238,  -12'd333,  12'd335,  12'd384,  -12'd51,  -12'd124,  12'd156,  12'd107,  12'd102,  12'd423,  -12'd27,  12'd323,  12'd320,  -12'd6,  12'd196,  
-12'd434,  12'd290,  12'd1,  12'd159,  12'd22,  12'd190,  -12'd43,  12'd173,  12'd55,  -12'd224,  -12'd3,  12'd119,  12'd182,  -12'd389,  12'd182,  12'd480,  
-12'd373,  -12'd137,  -12'd413,  12'd81,  -12'd97,  -12'd232,  -12'd286,  12'd133,  -12'd144,  12'd58,  -12'd49,  -12'd77,  12'd402,  -12'd201,  12'd184,  12'd201,  
12'd15,  -12'd379,  12'd215,  12'd43,  -12'd25,  12'd234,  12'd160,  -12'd30,  -12'd400,  -12'd197,  12'd172,  12'd68,  12'd193,  -12'd300,  -12'd379,  12'd181,  
-12'd47,  -12'd35,  12'd10,  12'd108,  12'd114,  12'd26,  -12'd16,  12'd325,  -12'd285,  12'd193,  -12'd21,  12'd232,  12'd52,  12'd39,  -12'd112,  12'd213,  
-12'd83,  -12'd364,  -12'd152,  12'd77,  -12'd231,  -12'd65,  12'd15,  12'd351,  -12'd393,  12'd7,  12'd313,  -12'd84,  12'd46,  -12'd224,  -12'd125,  -12'd101,  
-12'd262,  12'd87,  12'd104,  -12'd63,  -12'd26,  -12'd29,  -12'd73,  12'd69,  -12'd205,  12'd136,  12'd21,  -12'd175,  -12'd172,  12'd407,  -12'd273,  12'd321,  
-12'd116,  12'd440,  12'd205,  12'd177,  -12'd59,  -12'd138,  12'd315,  12'd128,  -12'd224,  -12'd52,  12'd20,  12'd358,  12'd159,  12'd171,  12'd119,  -12'd42,  
12'd10,  12'd386,  12'd126,  -12'd49,  12'd196,  -12'd122,  -12'd311,  12'd380,  -12'd401,  -12'd43,  -12'd77,  -12'd85,  -12'd238,  -12'd72,  12'd189,  12'd156,  
12'd101,  -12'd27,  -12'd142,  -12'd14,  -12'd425,  12'd60,  -12'd81,  -12'd416,  12'd313,  12'd65,  12'd124,  -12'd14,  -12'd311,  -12'd319,  -12'd380,  -12'd118,  
12'd227,  -12'd356,  -12'd92,  -12'd39,  -12'd92,  -12'd198,  12'd199,  12'd20,  -12'd5,  12'd49,  12'd243,  -12'd206,  12'd209,  -12'd138,  12'd22,  -12'd9,  
-12'd71,  -12'd189,  -12'd113,  12'd4,  -12'd17,  -12'd43,  12'd183,  -12'd40,  12'd234,  12'd161,  -12'd29,  -12'd161,  12'd177,  12'd245,  -12'd306,  12'd158,  
12'd384,  12'd190,  12'd224,  12'd77,  12'd147,  -12'd366,  12'd39,  12'd173,  -12'd20,  -12'd474,  -12'd222,  -12'd263,  -12'd355,  -12'd123,  12'd226,  -12'd272,  
-12'd126,  12'd102,  12'd273,  12'd124,  12'd486,  12'd201,  -12'd17,  -12'd46,  12'd217,  -12'd87,  -12'd288,  12'd187,  12'd259,  12'd149,  -12'd31,  -12'd133,  
-12'd102,  -12'd28,  -12'd207,  -12'd94,  12'd186,  12'd94,  12'd65,  12'd8,  12'd250,  12'd270,  12'd254,  12'd47,  12'd257,  -12'd269,  12'd42,  -12'd56,  
-12'd81,  -12'd161,  -12'd278,  12'd110,  -12'd85,  12'd139,  -12'd23,  -12'd1,  12'd250,  12'd226,  12'd36,  -12'd81,  12'd179,  12'd73,  12'd201,  -12'd180,  
12'd264,  12'd39,  -12'd68,  12'd165,  -12'd119,  12'd199,  -12'd132,  -12'd240,  12'd105,  12'd143,  -12'd117,  12'd30,  12'd183,  12'd613,  -12'd91,  12'd157,  
-12'd182,  -12'd111,  12'd295,  12'd249,  12'd25,  -12'd76,  12'd70,  -12'd289,  12'd181,  -12'd170,  12'd39,  12'd345,  12'd87,  -12'd67,  -12'd92,  -12'd155,  
-12'd123,  -12'd297,  12'd53,  12'd144,  12'd422,  -12'd157,  -12'd111,  12'd55,  12'd133,  12'd296,  -12'd29,  12'd253,  12'd271,  12'd79,  12'd44,  -12'd265,  
12'd14,  -12'd42,  12'd47,  -12'd230,  -12'd472,  -12'd128,  12'd285,  12'd14,  12'd71,  -12'd136,  12'd399,  -12'd319,  -12'd177,  12'd213,  -12'd109,  -12'd32,  
12'd12,  12'd100,  -12'd141,  12'd297,  -12'd166,  12'd269,  12'd459,  12'd440,  12'd135,  12'd110,  12'd334,  -12'd118,  12'd42,  12'd251,  12'd491,  12'd19,  
-12'd101,  -12'd280,  12'd220,  12'd179,  -12'd229,  -12'd313,  -12'd193,  -12'd194,  -12'd278,  -12'd227,  -12'd352,  -12'd181,  -12'd246,  12'd507,  12'd261,  12'd170,  
-12'd353,  12'd100,  -12'd104,  -12'd52,  12'd17,  -12'd71,  12'd151,  -12'd63,  -12'd18,  -12'd115,  -12'd62,  -12'd104,  12'd178,  -12'd147,  12'd134,  12'd165,  
12'd19,  12'd551,  -12'd43,  12'd88,  12'd384,  12'd283,  -12'd303,  -12'd168,  12'd85,  12'd330,  12'd63,  -12'd52,  -12'd114,  12'd196,  -12'd299,  12'd87,  

-12'd380,  -12'd14,  -12'd50,  -12'd57,  -12'd214,  12'd159,  12'd350,  12'd174,  -12'd285,  12'd69,  12'd126,  12'd51,  12'd124,  12'd269,  12'd60,  -12'd212,  
12'd354,  -12'd44,  12'd22,  -12'd32,  12'd202,  12'd172,  12'd321,  12'd176,  -12'd220,  12'd150,  12'd523,  12'd328,  -12'd66,  12'd116,  12'd101,  12'd113,  
12'd160,  12'd56,  -12'd39,  12'd291,  12'd377,  12'd132,  12'd221,  12'd38,  12'd132,  -12'd60,  12'd321,  12'd133,  -12'd38,  12'd261,  12'd241,  -12'd171,  
-12'd20,  12'd565,  12'd360,  -12'd29,  -12'd74,  12'd47,  -12'd256,  12'd93,  12'd79,  -12'd122,  -12'd134,  12'd235,  12'd138,  -12'd237,  -12'd286,  12'd353,  
-12'd53,  12'd92,  12'd174,  -12'd72,  -12'd32,  12'd1,  -12'd430,  12'd98,  12'd237,  12'd156,  12'd16,  12'd15,  -12'd31,  12'd200,  -12'd194,  -12'd113,  
12'd136,  -12'd94,  -12'd325,  -12'd11,  -12'd19,  -12'd408,  12'd7,  12'd5,  -12'd264,  -12'd58,  12'd302,  -12'd223,  12'd4,  12'd73,  -12'd240,  -12'd48,  
-12'd197,  -12'd48,  12'd505,  12'd216,  -12'd207,  12'd350,  12'd550,  -12'd210,  12'd20,  12'd80,  -12'd157,  -12'd25,  -12'd354,  12'd70,  12'd101,  -12'd210,  
-12'd361,  12'd470,  12'd11,  12'd35,  12'd317,  -12'd26,  12'd263,  -12'd144,  12'd264,  12'd142,  12'd284,  -12'd503,  -12'd87,  -12'd18,  -12'd142,  -12'd222,  
-12'd576,  -12'd17,  -12'd239,  -12'd244,  12'd364,  -12'd153,  -12'd512,  -12'd160,  -12'd70,  12'd390,  -12'd139,  -12'd168,  -12'd371,  -12'd197,  12'd63,  -12'd30,  
-12'd1035,  -12'd483,  12'd336,  -12'd324,  -12'd390,  12'd2,  -12'd311,  -12'd88,  -12'd211,  -12'd108,  -12'd18,  -12'd378,  -12'd493,  -12'd28,  12'd456,  12'd59,  
-12'd20,  -12'd281,  -12'd162,  -12'd142,  -12'd340,  -12'd209,  12'd644,  -12'd224,  12'd165,  -12'd229,  -12'd20,  12'd166,  -12'd202,  -12'd155,  12'd7,  12'd114,  
12'd348,  -12'd303,  12'd46,  12'd30,  -12'd350,  -12'd202,  -12'd347,  12'd94,  12'd34,  12'd29,  -12'd244,  -12'd230,  -12'd66,  -12'd118,  -12'd366,  -12'd99,  
-12'd424,  -12'd28,  -12'd12,  -12'd56,  12'd133,  -12'd416,  -12'd298,  12'd114,  12'd263,  12'd238,  -12'd426,  -12'd70,  -12'd408,  12'd85,  -12'd35,  -12'd139,  
-12'd121,  12'd235,  12'd142,  -12'd35,  -12'd220,  12'd101,  12'd47,  -12'd503,  12'd285,  -12'd224,  -12'd368,  12'd79,  -12'd214,  12'd296,  -12'd122,  -12'd456,  
-12'd158,  -12'd71,  12'd512,  12'd32,  -12'd148,  -12'd58,  -12'd39,  -12'd34,  12'd274,  12'd32,  -12'd385,  12'd599,  -12'd375,  12'd311,  12'd247,  -12'd558,  
12'd429,  12'd177,  12'd196,  -12'd88,  -12'd406,  12'd129,  12'd11,  12'd179,  12'd22,  12'd327,  -12'd406,  12'd25,  12'd371,  12'd176,  12'd99,  12'd32,  
-12'd83,  -12'd4,  12'd114,  -12'd149,  -12'd300,  12'd224,  12'd142,  12'd250,  12'd178,  -12'd60,  12'd230,  12'd202,  -12'd192,  12'd580,  12'd290,  12'd453,  
12'd116,  -12'd396,  12'd137,  12'd195,  -12'd182,  12'd150,  -12'd89,  12'd134,  -12'd118,  12'd63,  12'd86,  12'd164,  12'd27,  12'd130,  -12'd126,  12'd343,  
12'd24,  12'd200,  12'd288,  12'd307,  -12'd84,  -12'd25,  12'd78,  -12'd204,  12'd86,  -12'd136,  -12'd46,  12'd25,  12'd267,  12'd193,  12'd132,  -12'd132,  
12'd669,  -12'd2,  12'd243,  12'd404,  12'd154,  -12'd150,  12'd82,  -12'd23,  -12'd303,  12'd251,  12'd163,  12'd356,  12'd383,  -12'd373,  12'd40,  -12'd302,  
-12'd67,  -12'd61,  -12'd152,  12'd95,  -12'd149,  -12'd215,  -12'd11,  -12'd113,  -12'd255,  -12'd53,  -12'd205,  -12'd28,  -12'd109,  12'd17,  -12'd31,  12'd93,  
-12'd217,  12'd168,  -12'd87,  12'd298,  12'd5,  12'd31,  12'd212,  -12'd309,  -12'd86,  12'd34,  12'd83,  -12'd92,  -12'd43,  12'd412,  12'd208,  12'd38,  
-12'd18,  12'd239,  12'd235,  12'd104,  -12'd74,  12'd110,  12'd207,  12'd118,  12'd121,  12'd109,  -12'd5,  -12'd154,  -12'd77,  -12'd240,  -12'd179,  12'd54,  
-12'd73,  12'd403,  -12'd144,  -12'd82,  12'd16,  -12'd160,  -12'd251,  12'd59,  12'd32,  -12'd316,  -12'd0,  -12'd417,  12'd208,  -12'd236,  -12'd77,  12'd359,  
-12'd118,  12'd237,  -12'd434,  -12'd76,  12'd177,  -12'd159,  -12'd61,  12'd170,  -12'd224,  12'd10,  -12'd195,  -12'd81,  -12'd68,  -12'd65,  -12'd105,  12'd31,  

-12'd72,  12'd378,  -12'd128,  -12'd78,  12'd59,  -12'd26,  -12'd169,  -12'd50,  12'd137,  12'd56,  -12'd162,  -12'd83,  12'd356,  -12'd301,  12'd92,  12'd140,  
-12'd137,  -12'd91,  -12'd381,  12'd47,  12'd113,  12'd233,  -12'd247,  12'd69,  -12'd66,  -12'd176,  -12'd313,  12'd92,  12'd259,  -12'd84,  12'd285,  12'd223,  
-12'd136,  -12'd199,  12'd157,  12'd139,  -12'd138,  -12'd139,  12'd330,  12'd28,  -12'd365,  -12'd12,  12'd209,  -12'd81,  12'd177,  -12'd510,  12'd25,  12'd97,  
-12'd192,  -12'd147,  -12'd145,  -12'd108,  -12'd151,  12'd182,  12'd386,  -12'd279,  12'd189,  -12'd16,  12'd292,  12'd173,  -12'd357,  12'd235,  -12'd238,  12'd99,  
-12'd94,  12'd265,  -12'd240,  12'd12,  -12'd159,  -12'd121,  12'd259,  12'd10,  -12'd166,  -12'd206,  12'd9,  -12'd20,  -12'd295,  12'd32,  -12'd417,  12'd27,  
12'd107,  12'd50,  12'd12,  12'd346,  -12'd24,  -12'd89,  -12'd278,  12'd306,  -12'd218,  -12'd573,  12'd209,  12'd49,  -12'd187,  12'd185,  -12'd55,  12'd168,  
-12'd284,  12'd126,  12'd7,  -12'd82,  12'd60,  12'd294,  -12'd69,  -12'd33,  -12'd249,  12'd96,  12'd265,  -12'd29,  12'd263,  -12'd435,  12'd265,  12'd322,  
-12'd92,  12'd1,  -12'd336,  -12'd272,  12'd380,  -12'd243,  12'd74,  -12'd54,  12'd106,  -12'd132,  12'd300,  12'd28,  -12'd171,  -12'd212,  -12'd28,  12'd400,  
12'd66,  -12'd109,  -12'd166,  -12'd244,  -12'd151,  12'd172,  12'd248,  12'd92,  12'd218,  12'd215,  12'd65,  -12'd161,  -12'd15,  12'd148,  -12'd72,  -12'd131,  
12'd261,  12'd343,  12'd314,  12'd224,  12'd8,  -12'd150,  -12'd261,  12'd152,  -12'd26,  12'd326,  12'd39,  -12'd374,  12'd283,  12'd134,  -12'd91,  -12'd134,  
12'd242,  12'd9,  12'd166,  -12'd182,  -12'd343,  -12'd195,  -12'd243,  12'd135,  12'd156,  12'd58,  12'd189,  -12'd331,  12'd321,  12'd104,  12'd33,  -12'd106,  
-12'd87,  12'd168,  -12'd106,  12'd10,  12'd215,  -12'd32,  -12'd430,  -12'd11,  -12'd249,  12'd72,  12'd37,  12'd207,  12'd157,  -12'd192,  -12'd171,  12'd70,  
-12'd316,  -12'd218,  12'd343,  -12'd194,  -12'd41,  12'd290,  -12'd194,  -12'd26,  -12'd376,  -12'd77,  -12'd134,  12'd19,  12'd229,  -12'd12,  12'd233,  -12'd211,  
-12'd163,  -12'd244,  -12'd347,  12'd156,  12'd196,  12'd73,  12'd2,  -12'd403,  12'd41,  12'd243,  -12'd107,  -12'd141,  12'd106,  -12'd420,  12'd15,  12'd135,  
-12'd479,  -12'd230,  12'd234,  12'd201,  -12'd29,  -12'd13,  -12'd301,  -12'd2,  12'd209,  12'd581,  -12'd3,  12'd156,  -12'd244,  12'd339,  -12'd241,  -12'd240,  
-12'd448,  12'd101,  -12'd23,  12'd9,  -12'd49,  -12'd11,  -12'd217,  -12'd123,  12'd604,  -12'd16,  12'd248,  -12'd511,  -12'd248,  -12'd398,  -12'd207,  -12'd416,  
-12'd255,  -12'd135,  -12'd292,  -12'd160,  -12'd252,  12'd92,  -12'd209,  -12'd168,  -12'd129,  12'd412,  12'd334,  -12'd320,  12'd117,  -12'd329,  -12'd312,  -12'd223,  
-12'd22,  -12'd74,  12'd167,  -12'd80,  12'd93,  -12'd161,  -12'd123,  -12'd22,  -12'd138,  -12'd66,  12'd39,  -12'd81,  -12'd135,  -12'd276,  -12'd93,  12'd164,  
-12'd116,  -12'd3,  -12'd213,  12'd236,  12'd396,  12'd250,  -12'd340,  12'd27,  -12'd186,  -12'd263,  -12'd173,  12'd261,  12'd394,  -12'd277,  -12'd65,  12'd91,  
-12'd356,  -12'd67,  12'd72,  12'd299,  -12'd38,  12'd172,  12'd119,  -12'd113,  12'd167,  12'd214,  -12'd51,  12'd139,  12'd40,  12'd84,  -12'd252,  -12'd303,  
-12'd74,  -12'd90,  -12'd310,  12'd255,  12'd107,  12'd170,  12'd564,  -12'd220,  12'd303,  12'd94,  12'd442,  -12'd215,  -12'd114,  -12'd153,  -12'd32,  -12'd254,  
12'd311,  12'd42,  -12'd64,  -12'd48,  -12'd235,  -12'd329,  12'd17,  -12'd285,  12'd556,  12'd397,  -12'd44,  12'd221,  12'd162,  -12'd570,  -12'd110,  12'd19,  
12'd142,  12'd277,  -12'd170,  12'd225,  12'd3,  12'd19,  -12'd127,  -12'd28,  12'd383,  12'd501,  12'd217,  12'd307,  -12'd177,  12'd90,  -12'd201,  12'd265,  
12'd402,  12'd275,  -12'd261,  -12'd212,  12'd251,  12'd301,  -12'd118,  12'd190,  12'd175,  -12'd209,  -12'd26,  -12'd225,  12'd380,  12'd324,  -12'd60,  -12'd150,  
12'd100,  12'd81,  12'd374,  12'd101,  -12'd48,  12'd185,  -12'd154,  -12'd239,  12'd356,  12'd62,  -12'd95,  -12'd246,  -12'd54,  12'd265,  -12'd285,  12'd180,  

12'd436,  -12'd438,  -12'd242,  12'd28,  -12'd382,  12'd221,  12'd96,  -12'd136,  -12'd257,  12'd146,  12'd310,  12'd53,  -12'd189,  12'd211,  -12'd396,  -12'd185,  
-12'd101,  -12'd171,  -12'd32,  -12'd325,  -12'd278,  12'd89,  12'd62,  -12'd526,  12'd30,  -12'd60,  -12'd69,  12'd381,  -12'd80,  12'd125,  12'd82,  12'd35,  
12'd174,  12'd0,  -12'd43,  -12'd142,  12'd165,  -12'd133,  -12'd328,  12'd291,  12'd358,  -12'd75,  -12'd93,  12'd183,  12'd139,  -12'd93,  -12'd75,  12'd309,  
-12'd21,  12'd84,  -12'd104,  12'd130,  -12'd131,  -12'd41,  12'd79,  12'd110,  12'd184,  -12'd184,  -12'd385,  -12'd181,  -12'd299,  12'd124,  12'd164,  12'd189,  
-12'd292,  12'd81,  -12'd0,  12'd41,  12'd42,  -12'd67,  12'd269,  12'd12,  12'd143,  -12'd27,  -12'd310,  12'd89,  12'd0,  12'd179,  -12'd325,  -12'd230,  
12'd51,  -12'd76,  12'd106,  12'd174,  12'd95,  12'd195,  12'd439,  -12'd234,  12'd374,  -12'd147,  12'd100,  12'd360,  -12'd21,  12'd192,  -12'd234,  -12'd278,  
12'd65,  12'd141,  12'd80,  12'd167,  -12'd3,  -12'd52,  12'd234,  -12'd288,  12'd493,  12'd211,  -12'd479,  12'd60,  -12'd78,  12'd261,  12'd320,  12'd283,  
12'd341,  12'd283,  12'd38,  -12'd12,  12'd256,  -12'd65,  12'd315,  12'd45,  -12'd268,  -12'd145,  -12'd99,  12'd160,  -12'd177,  -12'd62,  12'd91,  -12'd3,  
-12'd242,  -12'd195,  12'd12,  12'd35,  12'd259,  -12'd162,  12'd6,  -12'd377,  12'd199,  -12'd118,  -12'd387,  12'd218,  -12'd5,  12'd191,  -12'd219,  12'd209,  
12'd408,  -12'd118,  -12'd338,  12'd322,  -12'd160,  -12'd329,  12'd271,  -12'd150,  12'd4,  -12'd362,  12'd185,  12'd127,  12'd116,  -12'd36,  12'd143,  12'd211,  
12'd184,  12'd111,  12'd502,  12'd43,  12'd130,  12'd78,  12'd258,  12'd206,  -12'd198,  12'd103,  -12'd478,  12'd374,  12'd78,  12'd134,  12'd35,  12'd309,  
12'd155,  12'd50,  12'd44,  12'd48,  12'd371,  -12'd27,  12'd55,  12'd186,  12'd101,  12'd76,  -12'd210,  12'd103,  12'd87,  12'd61,  -12'd249,  -12'd63,  
12'd176,  -12'd32,  -12'd72,  12'd118,  -12'd437,  12'd244,  12'd246,  12'd43,  -12'd276,  -12'd362,  -12'd160,  12'd107,  -12'd402,  -12'd182,  -12'd151,  12'd161,  
12'd181,  -12'd30,  -12'd289,  -12'd26,  -12'd318,  12'd181,  12'd21,  12'd28,  12'd56,  -12'd122,  12'd1,  12'd93,  12'd190,  12'd247,  -12'd92,  -12'd172,  
-12'd2,  -12'd4,  -12'd267,  -12'd2,  12'd303,  12'd233,  -12'd12,  -12'd154,  -12'd291,  -12'd94,  12'd15,  -12'd106,  12'd440,  -12'd13,  -12'd208,  12'd202,  
12'd236,  12'd114,  12'd347,  12'd31,  12'd194,  -12'd15,  12'd72,  12'd170,  -12'd317,  12'd195,  -12'd478,  12'd405,  12'd247,  12'd162,  12'd170,  12'd3,  
12'd174,  12'd300,  -12'd10,  -12'd306,  -12'd81,  12'd16,  12'd61,  -12'd0,  -12'd272,  12'd42,  -12'd240,  -12'd382,  12'd340,  12'd72,  -12'd53,  12'd233,  
12'd358,  -12'd10,  -12'd173,  -12'd116,  -12'd228,  -12'd258,  12'd27,  12'd288,  -12'd172,  -12'd113,  12'd8,  -12'd227,  -12'd361,  12'd180,  -12'd132,  12'd116,  
12'd17,  12'd25,  -12'd101,  -12'd230,  12'd308,  -12'd458,  12'd304,  -12'd39,  -12'd193,  -12'd15,  12'd27,  -12'd147,  -12'd313,  -12'd345,  12'd75,  12'd172,  
-12'd337,  -12'd230,  -12'd103,  12'd314,  -12'd122,  -12'd224,  -12'd123,  -12'd200,  12'd38,  -12'd153,  12'd156,  12'd39,  -12'd338,  -12'd80,  -12'd193,  12'd65,  
12'd254,  12'd41,  12'd48,  12'd330,  -12'd153,  12'd259,  -12'd259,  12'd85,  -12'd661,  12'd368,  -12'd266,  -12'd27,  -12'd141,  12'd505,  12'd55,  -12'd38,  
12'd134,  -12'd269,  12'd216,  -12'd89,  -12'd326,  -12'd261,  -12'd200,  12'd305,  12'd27,  12'd21,  -12'd251,  -12'd132,  12'd153,  12'd338,  -12'd196,  -12'd65,  
-12'd165,  12'd98,  12'd4,  12'd126,  -12'd4,  12'd45,  -12'd437,  12'd245,  -12'd121,  -12'd233,  -12'd274,  -12'd145,  12'd216,  12'd107,  12'd364,  -12'd202,  
12'd26,  -12'd163,  12'd162,  12'd150,  12'd276,  -12'd218,  -12'd134,  -12'd116,  -12'd408,  -12'd243,  12'd31,  -12'd249,  -12'd200,  -12'd272,  12'd248,  -12'd165,  
-12'd104,  -12'd100,  -12'd123,  12'd54,  12'd64,  12'd272,  12'd69,  12'd89,  -12'd267,  -12'd480,  12'd70,  12'd215,  -12'd42,  -12'd91,  12'd271,  -12'd107,  

-12'd366,  -12'd211,  12'd34,  -12'd155,  -12'd361,  -12'd109,  12'd279,  12'd136,  12'd206,  -12'd93,  -12'd325,  -12'd135,  -12'd530,  -12'd23,  -12'd123,  -12'd475,  
-12'd255,  12'd59,  -12'd408,  12'd261,  12'd18,  -12'd17,  12'd41,  12'd113,  12'd263,  -12'd220,  -12'd116,  -12'd180,  -12'd193,  -12'd16,  12'd234,  -12'd138,  
12'd86,  -12'd245,  12'd164,  -12'd207,  -12'd203,  -12'd99,  -12'd505,  -12'd112,  12'd235,  12'd37,  -12'd106,  -12'd116,  12'd56,  -12'd219,  -12'd167,  12'd45,  
-12'd316,  -12'd43,  -12'd119,  12'd77,  12'd189,  -12'd370,  -12'd120,  12'd288,  -12'd351,  12'd245,  -12'd266,  12'd6,  12'd383,  -12'd548,  12'd48,  12'd325,  
-12'd280,  -12'd546,  12'd156,  -12'd71,  12'd274,  12'd52,  -12'd11,  -12'd62,  12'd69,  -12'd350,  12'd10,  -12'd129,  -12'd10,  12'd358,  12'd243,  12'd67,  
-12'd106,  -12'd190,  -12'd391,  -12'd84,  12'd86,  -12'd238,  12'd81,  -12'd16,  -12'd41,  -12'd72,  -12'd69,  -12'd95,  -12'd138,  12'd5,  -12'd459,  -12'd239,  
-12'd118,  12'd50,  -12'd71,  -12'd170,  -12'd22,  -12'd215,  -12'd549,  -12'd153,  -12'd319,  12'd455,  12'd5,  12'd165,  -12'd334,  12'd167,  -12'd387,  12'd366,  
-12'd62,  -12'd112,  -12'd193,  -12'd318,  12'd167,  12'd259,  -12'd93,  12'd240,  12'd275,  12'd149,  -12'd204,  12'd396,  12'd56,  12'd13,  12'd352,  -12'd241,  
-12'd218,  -12'd475,  -12'd276,  12'd97,  -12'd186,  12'd194,  -12'd161,  -12'd57,  -12'd118,  -12'd122,  12'd83,  12'd12,  -12'd75,  -12'd257,  12'd33,  12'd240,  
-12'd47,  -12'd49,  12'd272,  12'd230,  12'd186,  12'd158,  12'd181,  12'd265,  -12'd352,  -12'd91,  12'd362,  12'd371,  12'd459,  -12'd287,  -12'd10,  12'd232,  
12'd131,  12'd51,  -12'd277,  12'd283,  12'd52,  12'd212,  -12'd26,  12'd55,  12'd262,  -12'd323,  -12'd617,  12'd17,  12'd231,  -12'd234,  -12'd41,  -12'd274,  
-12'd328,  12'd190,  12'd255,  -12'd250,  -12'd95,  12'd167,  12'd124,  -12'd339,  12'd231,  12'd90,  12'd75,  12'd136,  -12'd73,  -12'd182,  12'd217,  -12'd331,  
12'd138,  12'd102,  12'd180,  -12'd195,  12'd23,  -12'd124,  -12'd159,  -12'd477,  -12'd248,  12'd449,  12'd392,  12'd177,  -12'd20,  12'd3,  -12'd25,  12'd144,  
12'd200,  12'd20,  12'd254,  12'd19,  -12'd62,  -12'd281,  12'd91,  12'd370,  -12'd19,  12'd152,  12'd218,  -12'd185,  -12'd10,  12'd379,  -12'd296,  12'd208,  
-12'd96,  -12'd176,  -12'd518,  -12'd251,  12'd209,  -12'd119,  -12'd115,  -12'd2,  -12'd417,  -12'd89,  12'd44,  -12'd335,  12'd122,  12'd91,  12'd245,  12'd328,  
12'd265,  -12'd65,  12'd149,  12'd187,  12'd191,  12'd402,  -12'd312,  -12'd114,  12'd439,  -12'd56,  -12'd163,  -12'd199,  -12'd297,  -12'd40,  12'd232,  -12'd187,  
-12'd234,  12'd212,  12'd144,  -12'd3,  12'd96,  12'd171,  -12'd272,  -12'd231,  12'd466,  12'd159,  12'd110,  -12'd360,  -12'd164,  -12'd177,  -12'd12,  12'd72,  
12'd252,  -12'd116,  -12'd60,  12'd118,  12'd415,  -12'd18,  12'd118,  12'd208,  -12'd61,  -12'd150,  12'd30,  12'd132,  -12'd69,  -12'd9,  12'd18,  12'd205,  
-12'd215,  -12'd78,  -12'd128,  -12'd177,  12'd157,  -12'd278,  12'd356,  -12'd342,  12'd170,  12'd191,  -12'd13,  12'd73,  -12'd47,  12'd32,  12'd88,  -12'd177,  
-12'd221,  -12'd432,  -12'd60,  -12'd229,  -12'd460,  -12'd67,  -12'd220,  -12'd37,  -12'd404,  -12'd493,  -12'd310,  -12'd52,  -12'd384,  12'd51,  -12'd249,  -12'd248,  
-12'd85,  -12'd114,  12'd160,  12'd156,  12'd499,  12'd168,  -12'd64,  12'd167,  12'd86,  -12'd173,  12'd261,  -12'd91,  12'd318,  -12'd78,  -12'd55,  -12'd224,  
12'd14,  12'd7,  12'd175,  12'd64,  12'd285,  -12'd66,  -12'd280,  12'd41,  -12'd346,  -12'd232,  12'd15,  -12'd92,  12'd71,  -12'd496,  12'd159,  -12'd144,  
12'd198,  -12'd191,  12'd218,  12'd160,  -12'd442,  12'd319,  12'd188,  -12'd263,  -12'd144,  -12'd463,  12'd129,  -12'd9,  -12'd77,  -12'd98,  -12'd186,  -12'd130,  
-12'd26,  -12'd231,  12'd25,  12'd347,  -12'd328,  12'd346,  12'd283,  -12'd446,  12'd424,  -12'd618,  -12'd156,  12'd300,  -12'd440,  12'd102,  -12'd277,  -12'd180,  
12'd83,  -12'd94,  12'd805,  12'd66,  -12'd213,  12'd19,  -12'd19,  -12'd234,  12'd708,  12'd369,  -12'd21,  -12'd304,  -12'd333,  12'd303,  -12'd667,  -12'd332,  

12'd37,  12'd121,  -12'd335,  12'd144,  -12'd268,  12'd44,  12'd324,  12'd138,  12'd143,  12'd86,  -12'd178,  -12'd157,  12'd27,  12'd173,  12'd29,  12'd162,  
12'd188,  -12'd208,  -12'd179,  -12'd141,  -12'd32,  12'd5,  12'd273,  -12'd247,  12'd444,  12'd124,  -12'd383,  -12'd107,  12'd82,  12'd263,  12'd406,  -12'd17,  
-12'd237,  -12'd33,  12'd3,  -12'd286,  12'd18,  -12'd218,  12'd210,  -12'd144,  -12'd281,  12'd177,  12'd38,  12'd149,  -12'd115,  -12'd47,  -12'd240,  12'd171,  
-12'd127,  12'd188,  12'd140,  -12'd27,  -12'd93,  -12'd384,  12'd214,  -12'd139,  12'd208,  -12'd331,  12'd63,  12'd143,  12'd119,  -12'd6,  -12'd213,  12'd373,  
12'd113,  12'd519,  -12'd228,  12'd290,  12'd288,  12'd18,  12'd29,  12'd208,  -12'd188,  12'd51,  12'd67,  12'd44,  12'd51,  -12'd170,  12'd224,  12'd294,  
-12'd228,  12'd319,  12'd72,  12'd49,  12'd4,  -12'd233,  12'd222,  12'd97,  -12'd109,  12'd355,  -12'd104,  -12'd407,  12'd165,  12'd168,  12'd226,  -12'd92,  
-12'd108,  -12'd412,  -12'd7,  12'd91,  12'd220,  12'd79,  -12'd343,  12'd16,  -12'd558,  12'd327,  -12'd138,  -12'd154,  12'd113,  12'd604,  12'd289,  -12'd188,  
12'd97,  -12'd164,  -12'd13,  12'd343,  12'd161,  -12'd79,  12'd265,  12'd446,  -12'd210,  -12'd377,  -12'd166,  12'd250,  -12'd63,  -12'd159,  12'd314,  12'd137,  
12'd22,  -12'd240,  12'd156,  12'd11,  -12'd104,  12'd12,  12'd271,  12'd269,  12'd345,  -12'd479,  12'd359,  12'd117,  -12'd57,  -12'd380,  12'd0,  -12'd362,  
12'd553,  -12'd255,  -12'd475,  -12'd279,  12'd92,  12'd271,  12'd94,  12'd247,  -12'd183,  -12'd302,  12'd107,  -12'd366,  12'd225,  12'd72,  -12'd584,  12'd95,  
-12'd307,  12'd144,  -12'd510,  12'd215,  12'd418,  -12'd72,  -12'd212,  -12'd57,  -12'd17,  -12'd314,  -12'd231,  -12'd229,  12'd336,  -12'd391,  -12'd252,  -12'd294,  
-12'd175,  12'd316,  -12'd108,  12'd239,  12'd40,  12'd105,  -12'd448,  12'd118,  -12'd86,  12'd113,  -12'd24,  -12'd52,  -12'd190,  12'd397,  12'd191,  12'd214,  
12'd451,  12'd370,  -12'd142,  12'd155,  12'd120,  12'd171,  -12'd118,  -12'd10,  12'd32,  12'd298,  12'd127,  -12'd218,  12'd264,  -12'd352,  12'd104,  -12'd131,  
-12'd557,  -12'd423,  -12'd287,  -12'd375,  12'd22,  -12'd383,  -12'd33,  -12'd19,  -12'd6,  -12'd75,  -12'd391,  -12'd483,  12'd257,  -12'd242,  -12'd193,  12'd25,  
-12'd391,  -12'd166,  -12'd321,  -12'd115,  -12'd38,  12'd13,  -12'd283,  12'd111,  -12'd312,  12'd207,  12'd225,  -12'd40,  -12'd302,  12'd43,  -12'd139,  12'd405,  
-12'd215,  -12'd249,  -12'd283,  12'd164,  12'd96,  -12'd83,  -12'd340,  -12'd337,  12'd71,  12'd189,  -12'd502,  12'd168,  -12'd69,  12'd119,  -12'd12,  12'd164,  
12'd195,  12'd337,  12'd431,  12'd94,  12'd416,  -12'd106,  12'd247,  -12'd98,  -12'd198,  12'd264,  -12'd249,  -12'd17,  -12'd23,  12'd173,  -12'd212,  12'd51,  
12'd155,  12'd255,  12'd176,  -12'd167,  12'd144,  12'd64,  12'd26,  -12'd309,  -12'd384,  -12'd23,  -12'd431,  12'd221,  12'd119,  -12'd412,  12'd46,  12'd108,  
12'd27,  -12'd300,  -12'd181,  12'd20,  12'd363,  12'd260,  12'd50,  -12'd170,  12'd162,  -12'd102,  -12'd262,  12'd287,  12'd49,  12'd278,  -12'd182,  -12'd135,  
-12'd157,  -12'd2,  12'd685,  -12'd197,  -12'd337,  -12'd5,  -12'd106,  -12'd75,  12'd41,  -12'd418,  -12'd85,  12'd155,  12'd9,  12'd265,  -12'd586,  -12'd350,  
-12'd81,  -12'd60,  12'd45,  -12'd12,  12'd341,  -12'd10,  -12'd563,  12'd119,  12'd621,  -12'd274,  -12'd49,  -12'd46,  -12'd9,  -12'd545,  12'd9,  -12'd47,  
12'd25,  -12'd102,  -12'd115,  12'd162,  12'd294,  12'd184,  -12'd185,  -12'd3,  12'd159,  12'd4,  12'd194,  12'd147,  12'd59,  -12'd506,  -12'd304,  12'd264,  
12'd336,  12'd189,  -12'd6,  -12'd181,  12'd141,  12'd40,  -12'd170,  -12'd4,  12'd12,  12'd397,  12'd212,  12'd482,  12'd307,  -12'd248,  -12'd296,  -12'd319,  
12'd78,  12'd96,  12'd286,  -12'd58,  -12'd224,  12'd386,  12'd276,  12'd96,  12'd386,  12'd202,  12'd290,  12'd399,  12'd232,  12'd364,  -12'd137,  -12'd139,  
12'd47,  12'd76,  12'd129,  -12'd303,  12'd58,  12'd213,  12'd257,  12'd252,  12'd592,  -12'd598,  12'd80,  12'd161,  12'd271,  12'd482,  -12'd403,  -12'd9,  

-12'd186,  12'd43,  -12'd323,  -12'd396,  -12'd329,  -12'd218,  12'd166,  -12'd105,  -12'd103,  -12'd185,  12'd95,  -12'd10,  -12'd156,  -12'd292,  -12'd180,  -12'd17,  
-12'd86,  12'd319,  12'd84,  -12'd71,  -12'd206,  -12'd158,  -12'd77,  -12'd70,  12'd146,  12'd65,  -12'd166,  -12'd268,  12'd1,  12'd169,  12'd175,  12'd48,  
-12'd144,  12'd288,  12'd219,  12'd123,  -12'd284,  12'd148,  12'd175,  12'd264,  -12'd308,  12'd200,  -12'd252,  -12'd280,  12'd120,  -12'd473,  -12'd119,  12'd219,  
-12'd204,  -12'd313,  12'd239,  12'd57,  12'd126,  12'd146,  -12'd170,  12'd43,  -12'd255,  -12'd74,  -12'd168,  12'd2,  -12'd119,  12'd187,  12'd88,  -12'd27,  
-12'd271,  -12'd6,  -12'd269,  -12'd44,  -12'd126,  -12'd146,  12'd5,  -12'd25,  12'd66,  12'd136,  12'd184,  -12'd345,  -12'd327,  12'd226,  -12'd144,  -12'd155,  
-12'd264,  12'd256,  12'd163,  12'd107,  -12'd280,  -12'd222,  12'd56,  -12'd165,  -12'd49,  -12'd555,  12'd410,  12'd242,  -12'd257,  12'd122,  12'd191,  -12'd306,  
12'd497,  12'd238,  12'd234,  12'd236,  -12'd93,  -12'd213,  12'd218,  12'd50,  12'd133,  -12'd201,  -12'd382,  -12'd26,  -12'd120,  12'd150,  12'd107,  -12'd238,  
12'd118,  -12'd178,  -12'd78,  -12'd108,  12'd50,  -12'd212,  -12'd189,  12'd134,  -12'd127,  -12'd190,  -12'd245,  12'd11,  12'd12,  -12'd365,  12'd111,  -12'd72,  
12'd150,  12'd50,  12'd5,  12'd126,  -12'd102,  -12'd219,  12'd43,  -12'd134,  -12'd293,  -12'd220,  -12'd45,  -12'd102,  -12'd147,  12'd153,  12'd183,  12'd341,  
-12'd160,  12'd411,  12'd430,  -12'd23,  -12'd172,  12'd41,  12'd88,  12'd455,  -12'd87,  12'd30,  -12'd223,  12'd20,  12'd89,  12'd106,  -12'd293,  12'd181,  
12'd207,  12'd36,  12'd198,  -12'd237,  -12'd394,  -12'd391,  12'd552,  -12'd111,  12'd248,  -12'd64,  -12'd574,  -12'd8,  12'd46,  12'd494,  12'd106,  -12'd295,  
12'd79,  12'd230,  12'd155,  -12'd15,  12'd69,  -12'd270,  12'd72,  12'd323,  12'd213,  12'd150,  -12'd325,  -12'd132,  -12'd305,  12'd141,  -12'd104,  12'd182,  
12'd72,  12'd352,  12'd45,  -12'd210,  -12'd185,  12'd196,  -12'd382,  12'd186,  -12'd177,  -12'd87,  -12'd300,  -12'd447,  12'd151,  12'd145,  12'd97,  -12'd58,  
12'd155,  12'd503,  -12'd9,  -12'd42,  12'd371,  12'd50,  12'd63,  12'd7,  -12'd300,  12'd271,  12'd347,  -12'd16,  12'd108,  12'd245,  12'd220,  12'd57,  
12'd277,  -12'd163,  12'd316,  12'd299,  12'd300,  12'd291,  12'd177,  12'd370,  -12'd196,  -12'd248,  12'd109,  -12'd180,  12'd64,  -12'd148,  12'd116,  12'd146,  
-12'd487,  -12'd69,  12'd173,  12'd292,  12'd68,  12'd352,  12'd4,  12'd158,  -12'd518,  -12'd115,  -12'd143,  -12'd134,  -12'd79,  12'd249,  -12'd202,  -12'd227,  
-12'd270,  12'd104,  12'd141,  12'd163,  12'd109,  -12'd160,  -12'd385,  12'd120,  -12'd959,  12'd19,  12'd205,  -12'd105,  12'd16,  -12'd119,  -12'd82,  -12'd414,  
12'd56,  12'd155,  12'd59,  12'd105,  -12'd289,  -12'd32,  12'd8,  -12'd13,  -12'd564,  -12'd92,  12'd284,  12'd95,  -12'd339,  -12'd383,  12'd121,  -12'd226,  
-12'd109,  12'd35,  -12'd160,  -12'd93,  -12'd269,  12'd228,  12'd224,  12'd161,  12'd123,  -12'd426,  12'd305,  12'd310,  12'd143,  -12'd155,  -12'd73,  12'd42,  
-12'd111,  -12'd95,  12'd64,  -12'd125,  -12'd86,  12'd141,  12'd360,  12'd326,  12'd4,  -12'd549,  -12'd128,  -12'd324,  -12'd91,  12'd33,  -12'd185,  -12'd42,  
-12'd230,  12'd352,  -12'd96,  12'd242,  12'd340,  12'd173,  -12'd343,  12'd106,  12'd144,  12'd10,  12'd287,  -12'd38,  12'd19,  -12'd357,  -12'd48,  -12'd34,  
-12'd336,  12'd255,  -12'd98,  12'd346,  12'd244,  12'd40,  12'd262,  12'd164,  12'd409,  -12'd135,  12'd176,  -12'd2,  -12'd210,  -12'd387,  12'd9,  -12'd86,  
12'd180,  12'd11,  -12'd129,  12'd342,  12'd196,  -12'd204,  12'd413,  12'd127,  12'd430,  -12'd16,  -12'd85,  12'd20,  -12'd35,  -12'd40,  -12'd173,  -12'd180,  
12'd39,  -12'd18,  -12'd31,  12'd59,  -12'd39,  -12'd129,  -12'd146,  12'd154,  12'd169,  12'd299,  -12'd315,  12'd21,  12'd247,  12'd263,  12'd94,  -12'd242,  
-12'd115,  12'd24,  -12'd362,  -12'd622,  -12'd236,  12'd83,  -12'd323,  -12'd363,  -12'd98,  -12'd196,  12'd83,  -12'd122,  -12'd221,  12'd202,  -12'd386,  -12'd58,  

-12'd25,  12'd273,  -12'd392,  -12'd161,  -12'd280,  12'd92,  -12'd80,  -12'd40,  -12'd81,  12'd16,  12'd268,  -12'd200,  -12'd246,  -12'd85,  12'd37,  12'd91,  
12'd68,  12'd84,  -12'd61,  12'd23,  -12'd215,  12'd412,  12'd233,  -12'd233,  -12'd66,  -12'd337,  -12'd102,  12'd42,  -12'd291,  12'd36,  -12'd453,  12'd147,  
-12'd303,  -12'd322,  -12'd312,  -12'd240,  12'd215,  12'd62,  12'd134,  12'd182,  12'd131,  12'd228,  12'd114,  12'd300,  12'd8,  12'd96,  12'd321,  -12'd197,  
12'd93,  12'd112,  12'd217,  -12'd298,  -12'd172,  -12'd244,  -12'd84,  12'd164,  12'd313,  12'd169,  -12'd14,  -12'd9,  -12'd115,  12'd386,  -12'd112,  12'd163,  
-12'd92,  12'd275,  12'd83,  12'd196,  12'd186,  12'd51,  12'd321,  -12'd145,  12'd181,  12'd294,  12'd215,  12'd206,  -12'd146,  -12'd116,  -12'd4,  -12'd378,  
12'd145,  -12'd43,  12'd68,  12'd175,  -12'd231,  12'd47,  12'd220,  -12'd22,  12'd367,  12'd452,  -12'd70,  12'd194,  -12'd94,  -12'd23,  -12'd175,  -12'd312,  
12'd42,  12'd129,  12'd138,  -12'd228,  12'd14,  12'd225,  12'd423,  12'd48,  12'd263,  -12'd235,  -12'd25,  12'd122,  -12'd105,  12'd411,  -12'd40,  12'd273,  
-12'd29,  -12'd14,  12'd351,  -12'd252,  -12'd204,  -12'd180,  12'd5,  -12'd21,  12'd46,  12'd190,  12'd71,  -12'd85,  -12'd64,  12'd57,  12'd135,  -12'd207,  
12'd280,  12'd184,  12'd115,  12'd80,  -12'd86,  -12'd195,  -12'd352,  -12'd488,  -12'd52,  -12'd10,  -12'd200,  -12'd80,  -12'd326,  12'd288,  12'd84,  12'd58,  
-12'd10,  -12'd98,  -12'd339,  -12'd33,  -12'd369,  12'd307,  12'd0,  -12'd46,  12'd280,  -12'd260,  12'd166,  -12'd49,  12'd86,  12'd74,  12'd165,  -12'd218,  
12'd275,  -12'd136,  12'd146,  12'd208,  12'd135,  -12'd74,  12'd73,  -12'd1,  12'd53,  -12'd227,  -12'd351,  12'd154,  12'd494,  12'd124,  12'd35,  12'd181,  
12'd90,  12'd352,  12'd10,  12'd5,  12'd325,  12'd3,  12'd74,  12'd164,  -12'd27,  12'd98,  12'd379,  12'd320,  -12'd30,  12'd422,  -12'd116,  -12'd108,  
-12'd10,  12'd134,  -12'd70,  -12'd42,  -12'd83,  12'd190,  12'd6,  12'd257,  -12'd444,  -12'd206,  -12'd27,  12'd147,  -12'd60,  12'd89,  -12'd35,  -12'd101,  
12'd569,  12'd240,  12'd25,  12'd224,  -12'd42,  -12'd73,  12'd121,  12'd168,  -12'd249,  -12'd566,  -12'd37,  -12'd25,  12'd16,  12'd168,  12'd234,  -12'd288,  
12'd87,  -12'd3,  -12'd453,  -12'd275,  -12'd187,  12'd99,  -12'd68,  -12'd96,  12'd259,  -12'd254,  -12'd152,  -12'd153,  12'd250,  12'd120,  -12'd24,  12'd373,  
12'd44,  12'd202,  -12'd21,  -12'd154,  12'd444,  12'd136,  -12'd67,  12'd125,  -12'd321,  -12'd71,  12'd68,  -12'd10,  -12'd5,  12'd314,  -12'd2,  12'd315,  
-12'd84,  -12'd185,  -12'd160,  -12'd94,  12'd541,  -12'd424,  -12'd73,  12'd83,  -12'd90,  -12'd103,  -12'd43,  -12'd45,  12'd270,  -12'd191,  -12'd194,  -12'd14,  
12'd169,  12'd310,  -12'd331,  12'd4,  12'd27,  -12'd22,  12'd158,  -12'd101,  12'd248,  -12'd9,  -12'd423,  12'd43,  -12'd264,  12'd201,  -12'd293,  12'd298,  
12'd40,  -12'd75,  12'd51,  -12'd122,  -12'd160,  12'd114,  -12'd234,  12'd177,  -12'd189,  -12'd60,  -12'd293,  -12'd29,  12'd293,  12'd66,  -12'd263,  -12'd65,  
12'd0,  -12'd342,  -12'd170,  -12'd108,  -12'd242,  -12'd233,  12'd314,  -12'd294,  -12'd104,  -12'd427,  12'd128,  12'd234,  12'd281,  -12'd48,  12'd4,  12'd152,  
12'd110,  12'd320,  12'd358,  12'd53,  -12'd259,  12'd99,  -12'd363,  12'd203,  -12'd615,  -12'd47,  12'd182,  -12'd5,  12'd147,  -12'd244,  -12'd83,  -12'd53,  
-12'd327,  -12'd212,  12'd16,  -12'd334,  12'd237,  -12'd308,  12'd240,  12'd193,  12'd275,  -12'd446,  -12'd354,  12'd26,  12'd165,  12'd212,  -12'd383,  -12'd97,  
-12'd517,  -12'd90,  -12'd233,  -12'd204,  -12'd48,  12'd160,  -12'd87,  12'd210,  12'd165,  -12'd339,  -12'd144,  -12'd203,  -12'd103,  12'd460,  12'd78,  12'd87,  
-12'd319,  -12'd310,  12'd286,  -12'd56,  12'd94,  -12'd283,  12'd183,  -12'd82,  -12'd132,  -12'd100,  -12'd419,  -12'd187,  12'd44,  12'd366,  -12'd278,  12'd8,  
12'd11,  -12'd78,  -12'd374,  12'd20,  12'd99,  -12'd6,  12'd0,  12'd275,  -12'd466,  -12'd24,  -12'd239,  12'd74,  12'd173,  -12'd245,  12'd33,  -12'd119,  

12'd153,  12'd205,  12'd140,  12'd36,  -12'd201,  12'd34,  -12'd422,  -12'd2,  12'd188,  -12'd231,  -12'd306,  12'd275,  12'd218,  -12'd95,  -12'd201,  12'd190,  
12'd14,  -12'd45,  -12'd59,  12'd233,  -12'd46,  -12'd100,  -12'd304,  -12'd47,  -12'd50,  12'd184,  12'd261,  12'd74,  12'd253,  12'd609,  -12'd360,  -12'd398,  
-12'd308,  12'd303,  12'd133,  -12'd196,  -12'd216,  12'd7,  -12'd318,  -12'd231,  12'd347,  -12'd124,  -12'd163,  -12'd65,  -12'd203,  12'd292,  12'd145,  -12'd39,  
12'd14,  12'd60,  -12'd62,  12'd102,  -12'd231,  12'd70,  -12'd295,  12'd62,  -12'd123,  -12'd131,  -12'd336,  12'd14,  -12'd234,  12'd191,  12'd426,  12'd189,  
12'd330,  12'd95,  -12'd392,  12'd426,  12'd177,  -12'd130,  -12'd99,  12'd109,  12'd278,  12'd173,  12'd131,  12'd47,  12'd289,  12'd305,  12'd282,  12'd125,  
12'd209,  -12'd315,  12'd136,  12'd203,  -12'd427,  12'd297,  -12'd195,  12'd340,  -12'd57,  12'd62,  -12'd371,  12'd40,  -12'd24,  12'd173,  12'd80,  12'd48,  
-12'd121,  -12'd544,  12'd411,  -12'd113,  12'd114,  12'd155,  12'd242,  -12'd80,  -12'd129,  -12'd159,  12'd134,  -12'd226,  12'd3,  12'd240,  12'd352,  12'd111,  
12'd188,  -12'd19,  -12'd32,  -12'd47,  -12'd247,  12'd122,  12'd94,  -12'd310,  -12'd104,  12'd287,  -12'd272,  -12'd78,  -12'd308,  12'd470,  12'd164,  -12'd358,  
-12'd68,  12'd137,  -12'd43,  -12'd42,  12'd19,  -12'd182,  12'd21,  -12'd70,  12'd280,  -12'd101,  12'd70,  12'd282,  -12'd202,  -12'd347,  12'd1,  -12'd120,  
12'd210,  12'd281,  -12'd122,  -12'd108,  -12'd402,  12'd363,  -12'd125,  -12'd174,  12'd450,  12'd8,  12'd205,  12'd53,  12'd73,  12'd428,  -12'd267,  12'd474,  
-12'd15,  12'd61,  -12'd3,  12'd408,  -12'd239,  12'd153,  12'd9,  12'd203,  12'd76,  12'd238,  12'd366,  -12'd99,  12'd68,  -12'd169,  12'd65,  -12'd49,  
12'd82,  12'd306,  12'd0,  12'd149,  12'd171,  12'd121,  -12'd21,  12'd288,  -12'd110,  12'd288,  -12'd202,  -12'd131,  -12'd145,  12'd331,  -12'd23,  12'd249,  
-12'd301,  12'd16,  -12'd60,  -12'd400,  12'd322,  12'd152,  12'd184,  12'd6,  -12'd214,  -12'd67,  12'd176,  -12'd152,  -12'd151,  12'd110,  -12'd166,  12'd29,  
-12'd443,  12'd312,  -12'd87,  -12'd161,  12'd208,  -12'd256,  -12'd133,  -12'd57,  -12'd282,  -12'd28,  -12'd167,  12'd400,  -12'd453,  -12'd113,  12'd271,  12'd217,  
-12'd198,  12'd225,  12'd169,  12'd201,  12'd56,  12'd145,  12'd67,  12'd212,  12'd127,  -12'd38,  -12'd184,  -12'd124,  -12'd337,  -12'd11,  -12'd119,  -12'd39,  
-12'd118,  12'd271,  12'd260,  12'd27,  12'd19,  12'd184,  12'd180,  12'd336,  12'd75,  -12'd141,  -12'd5,  12'd162,  12'd240,  -12'd356,  12'd126,  -12'd32,  
12'd152,  12'd80,  12'd84,  -12'd202,  12'd380,  -12'd197,  -12'd89,  -12'd82,  -12'd133,  12'd206,  12'd13,  12'd69,  12'd72,  12'd32,  12'd349,  -12'd147,  
12'd108,  -12'd48,  -12'd205,  -12'd26,  12'd63,  12'd24,  -12'd237,  12'd123,  -12'd444,  -12'd247,  12'd419,  12'd67,  12'd198,  12'd293,  -12'd260,  -12'd71,  
12'd90,  12'd250,  12'd126,  12'd287,  12'd240,  12'd145,  12'd7,  12'd411,  12'd157,  -12'd120,  -12'd48,  12'd245,  12'd111,  12'd134,  -12'd24,  -12'd22,  
12'd501,  12'd56,  -12'd101,  12'd188,  -12'd172,  -12'd26,  -12'd336,  12'd181,  12'd236,  12'd121,  -12'd1,  -12'd103,  -12'd196,  12'd203,  12'd74,  -12'd66,  
-12'd327,  12'd135,  -12'd308,  -12'd176,  -12'd350,  12'd228,  12'd521,  12'd21,  12'd315,  -12'd188,  12'd8,  -12'd110,  -12'd285,  -12'd76,  -12'd16,  12'd274,  
-12'd256,  -12'd158,  -12'd93,  -12'd247,  12'd174,  12'd375,  12'd106,  12'd105,  12'd66,  12'd24,  12'd287,  12'd17,  12'd273,  -12'd331,  12'd421,  -12'd86,  
12'd242,  -12'd79,  -12'd476,  -12'd417,  12'd132,  -12'd19,  -12'd127,  12'd23,  12'd28,  12'd127,  12'd56,  12'd255,  12'd34,  12'd76,  -12'd314,  -12'd272,  
12'd567,  12'd470,  12'd35,  12'd103,  12'd302,  12'd29,  12'd17,  12'd39,  -12'd101,  12'd374,  12'd154,  12'd178,  -12'd5,  12'd304,  12'd311,  -12'd44,  
-12'd223,  12'd392,  -12'd142,  12'd246,  -12'd137,  12'd99,  12'd240,  12'd489,  12'd218,  -12'd359,  -12'd203,  12'd442,  -12'd76,  -12'd238,  12'd156,  12'd278,  

-12'd136,  12'd236,  -12'd182,  -12'd68,  12'd284,  12'd188,  -12'd66,  12'd110,  12'd122,  -12'd9,  -12'd360,  -12'd68,  12'd87,  12'd141,  -12'd299,  12'd315,  
12'd206,  12'd200,  -12'd308,  -12'd175,  12'd57,  12'd141,  12'd24,  12'd176,  -12'd402,  -12'd181,  -12'd208,  -12'd222,  12'd79,  12'd51,  -12'd204,  -12'd236,  
-12'd247,  12'd215,  -12'd63,  12'd290,  -12'd193,  -12'd29,  12'd119,  -12'd22,  12'd83,  -12'd14,  -12'd12,  -12'd92,  12'd33,  12'd312,  12'd230,  -12'd312,  
12'd262,  -12'd22,  -12'd276,  -12'd169,  -12'd114,  12'd58,  12'd192,  -12'd264,  12'd19,  12'd170,  12'd155,  -12'd362,  -12'd176,  12'd79,  12'd14,  -12'd19,  
12'd152,  -12'd187,  12'd346,  12'd86,  12'd188,  -12'd261,  -12'd99,  12'd53,  -12'd301,  12'd66,  -12'd256,  -12'd130,  -12'd19,  -12'd312,  -12'd73,  12'd239,  
12'd32,  -12'd114,  12'd252,  -12'd6,  -12'd144,  -12'd70,  12'd163,  -12'd199,  -12'd14,  -12'd126,  12'd17,  12'd51,  -12'd153,  -12'd113,  12'd130,  -12'd39,  
-12'd87,  -12'd13,  -12'd238,  12'd150,  12'd69,  -12'd11,  -12'd82,  -12'd86,  -12'd172,  12'd115,  12'd93,  12'd224,  -12'd272,  12'd327,  -12'd60,  -12'd156,  
12'd31,  -12'd96,  12'd23,  -12'd440,  12'd137,  -12'd7,  12'd39,  -12'd385,  12'd95,  -12'd7,  -12'd155,  12'd70,  -12'd286,  12'd120,  12'd71,  -12'd176,  
-12'd21,  -12'd22,  12'd128,  12'd44,  12'd40,  -12'd346,  -12'd141,  -12'd167,  -12'd7,  -12'd168,  12'd77,  12'd63,  -12'd7,  12'd119,  12'd42,  12'd27,  
12'd92,  -12'd207,  12'd131,  12'd153,  12'd108,  12'd89,  -12'd146,  12'd74,  12'd355,  12'd87,  12'd60,  12'd16,  -12'd25,  12'd212,  -12'd131,  -12'd267,  
-12'd52,  -12'd217,  -12'd155,  12'd37,  -12'd118,  12'd128,  12'd165,  -12'd424,  -12'd45,  12'd132,  -12'd71,  12'd3,  12'd140,  12'd173,  12'd270,  -12'd292,  
12'd6,  -12'd21,  -12'd322,  -12'd84,  -12'd214,  -12'd260,  12'd245,  -12'd219,  -12'd390,  -12'd47,  12'd64,  -12'd110,  -12'd156,  12'd14,  -12'd360,  -12'd123,  
-12'd85,  12'd236,  12'd225,  12'd12,  -12'd156,  -12'd74,  -12'd197,  12'd106,  -12'd273,  -12'd396,  -12'd50,  12'd124,  12'd80,  12'd76,  -12'd307,  12'd199,  
-12'd77,  -12'd348,  12'd5,  -12'd118,  12'd44,  -12'd15,  12'd261,  -12'd267,  -12'd196,  -12'd123,  -12'd354,  12'd49,  -12'd162,  12'd269,  -12'd287,  -12'd252,  
-12'd151,  -12'd370,  -12'd134,  12'd0,  -12'd193,  12'd174,  -12'd163,  12'd83,  -12'd52,  -12'd265,  12'd66,  -12'd340,  -12'd229,  -12'd126,  12'd281,  12'd46,  
-12'd22,  12'd150,  12'd300,  -12'd282,  -12'd100,  12'd285,  -12'd385,  -12'd26,  -12'd320,  -12'd278,  12'd171,  -12'd317,  12'd72,  12'd324,  12'd171,  -12'd53,  
-12'd269,  -12'd223,  12'd59,  -12'd233,  -12'd258,  12'd7,  12'd341,  -12'd116,  12'd124,  12'd139,  12'd71,  12'd62,  -12'd50,  12'd290,  -12'd83,  12'd38,  
-12'd81,  12'd119,  -12'd258,  -12'd269,  12'd47,  -12'd30,  -12'd278,  12'd51,  -12'd85,  -12'd6,  12'd166,  12'd210,  -12'd225,  -12'd204,  -12'd258,  -12'd107,  
-12'd366,  -12'd95,  -12'd211,  12'd114,  12'd52,  12'd240,  -12'd31,  -12'd25,  -12'd88,  12'd91,  12'd148,  -12'd67,  -12'd54,  12'd44,  -12'd48,  -12'd199,  
-12'd207,  -12'd281,  12'd120,  12'd26,  12'd200,  12'd66,  12'd38,  -12'd48,  12'd100,  -12'd126,  -12'd346,  12'd156,  -12'd124,  12'd21,  -12'd184,  12'd103,  
-12'd27,  -12'd83,  12'd129,  12'd360,  12'd117,  -12'd201,  12'd113,  12'd5,  -12'd27,  12'd212,  12'd29,  -12'd6,  12'd49,  -12'd220,  -12'd216,  -12'd120,  
-12'd237,  -12'd34,  12'd317,  -12'd56,  -12'd88,  -12'd11,  -12'd248,  12'd16,  -12'd205,  12'd52,  12'd252,  -12'd42,  12'd53,  -12'd16,  -12'd80,  12'd163,  
-12'd93,  -12'd55,  12'd19,  -12'd84,  12'd116,  12'd190,  -12'd243,  12'd30,  12'd157,  -12'd221,  -12'd187,  -12'd321,  -12'd124,  -12'd374,  -12'd346,  -12'd49,  
-12'd82,  12'd339,  -12'd192,  12'd32,  -12'd87,  -12'd125,  12'd3,  12'd21,  12'd155,  12'd184,  -12'd227,  -12'd136,  -12'd424,  -12'd79,  -12'd190,  -12'd403,  
-12'd305,  12'd78,  -12'd117,  -12'd106,  -12'd340,  12'd142,  -12'd282,  12'd214,  -12'd158,  12'd267,  -12'd122,  -12'd231,  12'd6,  -12'd93,  -12'd384,  12'd53,  

-12'd140,  -12'd62,  12'd285,  -12'd268,  -12'd235,  12'd225,  12'd1,  -12'd283,  -12'd149,  12'd64,  12'd113,  -12'd101,  12'd37,  12'd278,  -12'd266,  -12'd192,  
-12'd46,  12'd45,  12'd221,  12'd128,  -12'd104,  -12'd17,  12'd171,  12'd133,  12'd142,  -12'd198,  -12'd18,  12'd317,  12'd127,  12'd269,  -12'd96,  -12'd44,  
12'd268,  12'd82,  12'd158,  12'd110,  12'd24,  12'd58,  12'd153,  -12'd19,  12'd68,  -12'd194,  -12'd66,  -12'd186,  12'd303,  -12'd64,  -12'd162,  12'd61,  
12'd364,  -12'd40,  -12'd316,  -12'd18,  -12'd233,  12'd73,  12'd315,  12'd134,  -12'd60,  -12'd322,  12'd38,  -12'd70,  12'd197,  -12'd616,  -12'd210,  12'd311,  
12'd258,  12'd426,  -12'd187,  12'd287,  12'd23,  -12'd77,  12'd305,  -12'd105,  12'd115,  12'd86,  -12'd12,  12'd267,  12'd283,  12'd338,  12'd57,  12'd614,  
12'd96,  12'd78,  12'd195,  -12'd29,  -12'd179,  12'd237,  -12'd72,  -12'd163,  -12'd81,  12'd87,  -12'd134,  12'd355,  12'd173,  12'd92,  -12'd162,  12'd353,  
-12'd161,  12'd173,  12'd156,  12'd286,  -12'd332,  12'd166,  12'd76,  12'd148,  12'd245,  -12'd361,  -12'd65,  12'd50,  -12'd207,  -12'd226,  -12'd126,  -12'd71,  
-12'd200,  12'd124,  -12'd182,  12'd37,  12'd348,  -12'd2,  -12'd130,  12'd334,  -12'd6,  12'd79,  -12'd237,  -12'd32,  12'd383,  -12'd132,  -12'd376,  -12'd85,  
12'd67,  12'd92,  -12'd403,  12'd172,  12'd167,  -12'd115,  -12'd372,  12'd99,  12'd83,  12'd379,  12'd370,  -12'd76,  12'd143,  -12'd549,  12'd367,  12'd243,  
-12'd50,  -12'd537,  -12'd196,  12'd462,  12'd401,  12'd236,  -12'd118,  -12'd108,  12'd22,  -12'd149,  12'd193,  12'd42,  12'd231,  12'd163,  12'd155,  12'd257,  
-12'd214,  12'd76,  -12'd82,  -12'd130,  -12'd445,  -12'd361,  12'd325,  12'd121,  12'd86,  12'd58,  -12'd498,  12'd48,  -12'd183,  12'd59,  12'd470,  12'd208,  
-12'd329,  12'd109,  -12'd105,  -12'd143,  -12'd53,  -12'd30,  12'd115,  12'd242,  12'd8,  12'd64,  -12'd180,  -12'd46,  -12'd448,  -12'd42,  12'd220,  -12'd281,  
-12'd227,  -12'd65,  12'd420,  12'd416,  -12'd251,  -12'd180,  12'd3,  -12'd17,  12'd180,  12'd362,  -12'd313,  -12'd180,  -12'd161,  12'd106,  12'd263,  -12'd66,  
-12'd112,  12'd89,  -12'd524,  -12'd107,  12'd265,  12'd76,  12'd223,  12'd67,  -12'd190,  12'd24,  -12'd96,  -12'd167,  12'd431,  -12'd317,  12'd233,  12'd331,  
-12'd618,  -12'd248,  12'd3,  -12'd82,  12'd258,  -12'd323,  -12'd299,  -12'd29,  12'd269,  12'd74,  12'd173,  -12'd193,  -12'd440,  -12'd152,  -12'd18,  12'd288,  
-12'd227,  12'd272,  12'd80,  12'd343,  -12'd92,  -12'd147,  -12'd124,  -12'd45,  -12'd165,  12'd34,  -12'd683,  -12'd41,  12'd52,  -12'd25,  12'd159,  12'd64,  
-12'd143,  -12'd251,  12'd177,  12'd8,  12'd167,  12'd281,  12'd13,  -12'd87,  -12'd574,  12'd165,  -12'd388,  -12'd208,  12'd378,  12'd10,  12'd113,  -12'd149,  
-12'd262,  12'd166,  12'd183,  -12'd119,  12'd263,  -12'd38,  -12'd192,  -12'd142,  -12'd258,  12'd146,  12'd340,  12'd376,  12'd89,  12'd480,  -12'd337,  12'd128,  
-12'd165,  -12'd189,  12'd230,  12'd145,  12'd112,  -12'd41,  12'd182,  -12'd241,  -12'd77,  -12'd52,  12'd519,  -12'd179,  -12'd63,  -12'd213,  12'd58,  12'd114,  
12'd38,  12'd320,  12'd27,  -12'd96,  12'd231,  12'd136,  12'd140,  12'd8,  12'd169,  -12'd146,  -12'd154,  12'd132,  -12'd10,  12'd116,  12'd40,  12'd35,  
-12'd146,  12'd205,  -12'd453,  -12'd18,  -12'd169,  -12'd79,  12'd135,  12'd74,  12'd312,  12'd105,  -12'd335,  -12'd53,  -12'd80,  12'd12,  -12'd168,  -12'd272,  
12'd146,  12'd179,  12'd155,  -12'd92,  -12'd23,  -12'd150,  12'd142,  12'd101,  12'd15,  -12'd284,  -12'd198,  12'd462,  -12'd168,  -12'd75,  12'd148,  12'd69,  
-12'd352,  12'd238,  -12'd330,  -12'd118,  -12'd306,  -12'd245,  12'd370,  -12'd19,  12'd71,  12'd186,  -12'd111,  -12'd112,  12'd145,  12'd117,  12'd126,  -12'd4,  
12'd101,  -12'd9,  12'd16,  -12'd138,  -12'd174,  -12'd282,  12'd45,  12'd229,  12'd161,  -12'd255,  12'd240,  12'd99,  -12'd301,  12'd304,  -12'd49,  -12'd103,  
12'd349,  -12'd149,  -12'd403,  -12'd123,  12'd9,  12'd78,  12'd367,  12'd187,  -12'd159,  -12'd381,  -12'd4,  -12'd202,  -12'd206,  12'd491,  -12'd36,  -12'd371,  

-12'd319,  -12'd241,  -12'd417,  -12'd136,  -12'd110,  -12'd171,  12'd680,  -12'd329,  12'd38,  12'd235,  -12'd95,  -12'd236,  -12'd142,  -12'd209,  -12'd310,  -12'd274,  
12'd78,  -12'd279,  12'd41,  12'd38,  -12'd118,  12'd3,  12'd59,  12'd61,  12'd366,  12'd168,  -12'd64,  -12'd170,  -12'd118,  12'd200,  -12'd437,  12'd15,  
12'd220,  12'd69,  -12'd220,  -12'd413,  12'd91,  -12'd38,  -12'd238,  -12'd201,  12'd87,  -12'd217,  12'd113,  -12'd328,  12'd183,  -12'd113,  -12'd8,  12'd187,  
12'd233,  12'd273,  12'd116,  12'd161,  12'd222,  12'd105,  -12'd240,  -12'd26,  12'd102,  12'd310,  12'd34,  12'd60,  -12'd131,  -12'd103,  12'd349,  -12'd13,  
-12'd507,  -12'd86,  12'd385,  12'd97,  12'd58,  12'd26,  -12'd47,  -12'd16,  -12'd278,  12'd381,  -12'd2,  -12'd18,  -12'd30,  -12'd130,  12'd145,  -12'd176,  
-12'd203,  12'd24,  12'd335,  12'd89,  -12'd266,  12'd105,  12'd72,  -12'd121,  -12'd117,  -12'd180,  12'd51,  -12'd55,  -12'd296,  -12'd224,  -12'd15,  -12'd56,  
12'd219,  12'd140,  -12'd146,  12'd439,  -12'd364,  12'd365,  -12'd322,  -12'd431,  12'd220,  -12'd42,  12'd108,  -12'd116,  12'd7,  -12'd360,  -12'd380,  -12'd99,  
-12'd9,  -12'd91,  12'd42,  12'd88,  12'd137,  -12'd140,  12'd72,  -12'd288,  -12'd50,  -12'd148,  12'd351,  -12'd103,  12'd218,  -12'd180,  -12'd239,  12'd406,  
-12'd288,  12'd259,  12'd97,  12'd160,  12'd141,  -12'd167,  12'd49,  12'd94,  -12'd79,  12'd103,  12'd43,  -12'd298,  -12'd115,  12'd210,  -12'd153,  12'd98,  
-12'd25,  -12'd79,  12'd401,  12'd128,  12'd108,  12'd295,  -12'd139,  12'd136,  -12'd96,  12'd161,  -12'd354,  12'd310,  -12'd207,  12'd101,  -12'd45,  -12'd390,  
12'd197,  12'd285,  -12'd192,  12'd298,  -12'd742,  -12'd336,  12'd169,  12'd23,  12'd3,  12'd51,  -12'd409,  12'd117,  12'd19,  -12'd205,  -12'd56,  -12'd9,  
12'd127,  12'd80,  12'd145,  -12'd64,  -12'd255,  -12'd106,  12'd170,  12'd129,  12'd618,  -12'd215,  12'd229,  -12'd228,  12'd46,  12'd286,  -12'd98,  12'd165,  
-12'd272,  12'd198,  -12'd40,  12'd197,  12'd456,  -12'd145,  12'd252,  12'd60,  12'd133,  12'd24,  12'd6,  12'd69,  12'd41,  -12'd26,  -12'd297,  -12'd153,  
12'd336,  -12'd106,  -12'd128,  -12'd79,  12'd130,  -12'd260,  -12'd100,  12'd261,  -12'd445,  -12'd45,  12'd128,  12'd184,  -12'd197,  12'd197,  12'd326,  -12'd292,  
12'd51,  12'd70,  12'd327,  12'd117,  12'd77,  12'd78,  -12'd91,  12'd161,  12'd390,  12'd91,  12'd69,  12'd51,  12'd328,  12'd193,  12'd289,  12'd115,  
-12'd17,  -12'd135,  12'd193,  12'd9,  -12'd239,  -12'd31,  12'd191,  12'd129,  12'd50,  -12'd91,  -12'd71,  12'd168,  12'd56,  12'd309,  12'd322,  -12'd239,  
12'd54,  12'd115,  12'd105,  12'd244,  -12'd202,  12'd60,  12'd99,  12'd19,  12'd272,  -12'd221,  12'd263,  -12'd47,  -12'd235,  -12'd130,  -12'd163,  -12'd271,  
-12'd260,  -12'd324,  -12'd282,  -12'd177,  -12'd10,  12'd337,  12'd208,  -12'd330,  -12'd52,  12'd180,  12'd448,  -12'd140,  -12'd122,  -12'd242,  -12'd80,  12'd206,  
-12'd243,  12'd295,  -12'd191,  -12'd235,  12'd20,  12'd281,  12'd64,  -12'd47,  -12'd126,  12'd338,  12'd67,  -12'd107,  12'd383,  12'd66,  -12'd75,  12'd5,  
12'd66,  -12'd95,  12'd88,  12'd19,  12'd238,  12'd320,  -12'd308,  12'd201,  12'd79,  12'd203,  12'd34,  12'd141,  12'd211,  -12'd300,  12'd293,  12'd555,  
-12'd112,  -12'd338,  12'd299,  12'd93,  12'd254,  -12'd85,  -12'd433,  12'd292,  -12'd7,  -12'd158,  12'd10,  -12'd6,  -12'd108,  12'd402,  12'd376,  -12'd48,  
-12'd481,  -12'd225,  -12'd57,  12'd144,  12'd8,  12'd177,  -12'd50,  12'd293,  -12'd152,  -12'd182,  12'd102,  -12'd26,  12'd129,  -12'd199,  12'd4,  -12'd254,  
-12'd188,  -12'd712,  -12'd150,  12'd119,  12'd68,  12'd192,  -12'd280,  -12'd209,  -12'd319,  -12'd39,  12'd188,  -12'd202,  12'd37,  -12'd307,  -12'd65,  12'd313,  
-12'd107,  12'd64,  12'd61,  -12'd309,  12'd225,  -12'd259,  12'd62,  12'd47,  12'd37,  12'd448,  12'd145,  12'd87,  -12'd126,  -12'd307,  12'd126,  -12'd169,  
-12'd380,  12'd66,  -12'd314,  -12'd324,  12'd254,  -12'd366,  -12'd231,  -12'd108,  12'd324,  12'd565,  -12'd85,  12'd97,  12'd229,  -12'd527,  12'd4,  -12'd179,  

-12'd309,  -12'd241,  12'd69,  -12'd159,  -12'd357,  12'd71,  -12'd438,  -12'd112,  -12'd269,  -12'd132,  -12'd195,  -12'd241,  12'd111,  12'd354,  12'd161,  12'd56,  
12'd3,  -12'd31,  12'd2,  -12'd227,  12'd0,  12'd53,  -12'd49,  12'd217,  -12'd269,  12'd436,  -12'd92,  -12'd144,  12'd309,  -12'd99,  -12'd356,  12'd180,  
-12'd161,  -12'd312,  12'd9,  -12'd222,  12'd37,  12'd252,  -12'd45,  12'd288,  12'd120,  -12'd96,  -12'd123,  -12'd8,  12'd390,  -12'd150,  12'd209,  -12'd153,  
-12'd127,  12'd437,  12'd39,  12'd112,  12'd35,  -12'd71,  -12'd397,  -12'd81,  -12'd102,  -12'd242,  12'd209,  -12'd35,  -12'd59,  -12'd518,  12'd417,  -12'd373,  
12'd429,  -12'd19,  -12'd16,  12'd499,  -12'd39,  -12'd44,  -12'd5,  -12'd90,  -12'd184,  -12'd61,  12'd250,  12'd185,  -12'd202,  -12'd127,  12'd293,  -12'd186,  
-12'd271,  -12'd168,  12'd34,  -12'd449,  -12'd164,  12'd163,  12'd69,  -12'd304,  12'd128,  -12'd189,  -12'd255,  -12'd67,  12'd11,  -12'd146,  12'd202,  12'd318,  
12'd378,  -12'd136,  12'd54,  12'd219,  -12'd138,  -12'd156,  12'd26,  12'd15,  -12'd242,  -12'd34,  -12'd1,  -12'd108,  12'd169,  12'd64,  12'd9,  12'd52,  
12'd556,  12'd160,  12'd53,  12'd33,  12'd4,  12'd164,  12'd703,  12'd16,  12'd69,  -12'd225,  -12'd436,  -12'd212,  -12'd91,  -12'd20,  12'd191,  -12'd497,  
12'd293,  12'd346,  12'd224,  12'd151,  12'd393,  12'd4,  -12'd35,  -12'd170,  12'd472,  12'd243,  12'd223,  12'd383,  -12'd78,  12'd365,  12'd374,  -12'd46,  
12'd42,  -12'd235,  -12'd40,  -12'd84,  -12'd196,  12'd135,  12'd171,  12'd213,  12'd440,  -12'd31,  12'd192,  12'd421,  -12'd120,  12'd147,  12'd22,  -12'd264,  
-12'd429,  -12'd74,  -12'd96,  12'd48,  -12'd506,  12'd108,  12'd101,  -12'd192,  -12'd275,  -12'd381,  -12'd155,  12'd50,  -12'd202,  12'd432,  12'd218,  -12'd48,  
12'd548,  12'd114,  -12'd35,  -12'd188,  -12'd266,  -12'd46,  -12'd17,  -12'd187,  -12'd50,  -12'd101,  -12'd23,  12'd388,  12'd62,  12'd81,  -12'd306,  12'd152,  
12'd192,  12'd407,  12'd187,  -12'd154,  12'd249,  12'd12,  12'd461,  -12'd22,  12'd108,  12'd49,  -12'd129,  12'd165,  12'd70,  12'd187,  12'd65,  -12'd71,  
12'd223,  12'd235,  12'd138,  -12'd124,  -12'd127,  12'd188,  -12'd75,  12'd13,  -12'd76,  -12'd405,  12'd376,  12'd177,  -12'd175,  -12'd51,  12'd259,  12'd176,  
12'd114,  12'd221,  -12'd75,  -12'd105,  -12'd152,  -12'd28,  -12'd48,  -12'd0,  12'd511,  -12'd145,  12'd225,  -12'd167,  -12'd44,  12'd365,  -12'd14,  -12'd315,  
12'd45,  -12'd121,  -12'd24,  12'd53,  -12'd147,  -12'd176,  12'd292,  -12'd258,  -12'd314,  -12'd141,  -12'd28,  12'd287,  12'd121,  -12'd26,  12'd115,  -12'd17,  
12'd425,  12'd267,  12'd127,  -12'd83,  -12'd152,  -12'd254,  12'd170,  12'd42,  -12'd342,  -12'd325,  -12'd133,  -12'd21,  12'd215,  -12'd68,  -12'd290,  12'd47,  
12'd209,  12'd110,  -12'd245,  12'd20,  -12'd330,  -12'd173,  12'd233,  -12'd110,  -12'd353,  -12'd192,  12'd389,  -12'd96,  -12'd80,  12'd352,  -12'd349,  -12'd235,  
12'd147,  12'd154,  12'd339,  -12'd48,  -12'd314,  12'd164,  12'd242,  12'd75,  -12'd114,  -12'd380,  12'd342,  -12'd0,  12'd75,  -12'd272,  12'd23,  12'd137,  
-12'd229,  -12'd184,  -12'd434,  -12'd486,  -12'd88,  -12'd425,  12'd161,  12'd78,  -12'd407,  -12'd802,  -12'd55,  -12'd452,  12'd148,  12'd90,  -12'd544,  -12'd38,  
-12'd168,  12'd95,  -12'd68,  -12'd69,  -12'd407,  -12'd18,  -12'd85,  12'd223,  -12'd244,  12'd161,  12'd268,  12'd190,  -12'd2,  12'd269,  12'd210,  -12'd32,  
12'd255,  -12'd123,  12'd418,  12'd79,  -12'd107,  -12'd76,  12'd176,  -12'd1,  -12'd292,  12'd137,  -12'd34,  -12'd247,  12'd109,  12'd158,  12'd96,  12'd176,  
-12'd276,  12'd281,  12'd58,  -12'd291,  12'd78,  -12'd565,  12'd322,  -12'd75,  -12'd183,  12'd519,  -12'd155,  -12'd343,  -12'd51,  12'd390,  -12'd253,  -12'd230,  
-12'd490,  -12'd487,  12'd31,  -12'd809,  -12'd208,  -12'd368,  12'd34,  -12'd27,  12'd6,  -12'd215,  -12'd322,  -12'd524,  -12'd273,  -12'd13,  -12'd342,  -12'd194,  
12'd53,  -12'd335,  -12'd423,  -12'd579,  -12'd541,  -12'd390,  -12'd307,  -12'd190,  -12'd325,  -12'd629,  -12'd211,  -12'd604,  -12'd722,  -12'd186,  -12'd353,  -12'd622,  

-12'd57,  12'd140,  12'd230,  12'd91,  -12'd191,  -12'd149,  -12'd34,  -12'd111,  12'd168,  -12'd62,  12'd65,  -12'd97,  12'd188,  12'd100,  -12'd138,  12'd291,  
12'd74,  12'd425,  12'd641,  12'd114,  12'd105,  -12'd161,  12'd245,  12'd86,  12'd281,  -12'd104,  12'd251,  12'd135,  12'd77,  12'd16,  -12'd168,  -12'd89,  
-12'd129,  12'd45,  12'd349,  -12'd58,  12'd230,  12'd378,  12'd388,  12'd138,  -12'd58,  -12'd593,  -12'd84,  12'd270,  -12'd131,  12'd776,  12'd214,  -12'd12,  
12'd267,  12'd8,  12'd31,  12'd102,  12'd240,  -12'd185,  -12'd161,  12'd247,  12'd124,  12'd373,  12'd168,  12'd199,  -12'd280,  12'd295,  12'd46,  12'd276,  
-12'd408,  -12'd183,  -12'd1,  12'd273,  -12'd650,  -12'd106,  -12'd183,  12'd196,  12'd32,  12'd259,  -12'd236,  12'd190,  -12'd324,  -12'd270,  12'd47,  -12'd250,  
-12'd168,  12'd444,  12'd254,  12'd97,  12'd203,  -12'd155,  12'd248,  -12'd35,  -12'd409,  -12'd268,  12'd37,  -12'd307,  -12'd246,  12'd292,  -12'd118,  -12'd149,  
12'd165,  -12'd99,  12'd76,  -12'd281,  12'd4,  12'd17,  12'd180,  -12'd284,  12'd8,  12'd128,  12'd560,  12'd19,  12'd273,  12'd446,  12'd86,  12'd55,  
-12'd169,  -12'd44,  12'd73,  12'd87,  -12'd223,  12'd190,  12'd84,  -12'd419,  12'd12,  -12'd113,  12'd108,  12'd7,  12'd235,  12'd123,  -12'd125,  12'd304,  
-12'd128,  12'd501,  -12'd269,  12'd136,  12'd501,  12'd22,  -12'd344,  -12'd62,  -12'd96,  12'd101,  -12'd0,  12'd127,  -12'd260,  -12'd244,  12'd79,  -12'd335,  
12'd222,  -12'd497,  12'd103,  -12'd13,  12'd140,  -12'd80,  12'd5,  -12'd264,  -12'd36,  12'd354,  -12'd38,  12'd7,  -12'd270,  12'd99,  12'd143,  -12'd167,  
12'd145,  12'd180,  12'd75,  -12'd439,  -12'd491,  -12'd486,  12'd540,  -12'd321,  -12'd453,  -12'd298,  12'd369,  12'd182,  -12'd518,  12'd312,  12'd149,  12'd130,  
12'd181,  -12'd93,  12'd345,  -12'd281,  -12'd228,  12'd63,  12'd266,  -12'd56,  12'd20,  -12'd75,  -12'd99,  -12'd108,  -12'd371,  12'd21,  -12'd154,  -12'd147,  
-12'd92,  12'd338,  -12'd198,  -12'd554,  12'd244,  -12'd314,  12'd88,  12'd145,  12'd331,  -12'd27,  -12'd179,  -12'd93,  -12'd247,  12'd75,  12'd190,  -12'd20,  
-12'd183,  12'd432,  -12'd87,  12'd170,  -12'd48,  -12'd227,  12'd287,  12'd141,  -12'd155,  -12'd243,  12'd67,  -12'd118,  -12'd179,  12'd86,  12'd96,  -12'd154,  
-12'd406,  12'd78,  12'd57,  -12'd237,  -12'd205,  -12'd227,  12'd117,  -12'd102,  12'd29,  -12'd361,  -12'd313,  -12'd7,  -12'd338,  -12'd185,  12'd181,  12'd153,  
12'd1,  -12'd174,  12'd249,  -12'd177,  -12'd196,  12'd227,  12'd112,  12'd165,  -12'd210,  12'd98,  12'd2,  -12'd107,  -12'd174,  12'd351,  -12'd159,  -12'd124,  
12'd185,  -12'd62,  12'd127,  -12'd513,  -12'd198,  -12'd0,  -12'd162,  -12'd128,  12'd145,  -12'd89,  -12'd134,  12'd16,  -12'd479,  12'd76,  -12'd185,  -12'd282,  
12'd347,  -12'd194,  12'd262,  12'd254,  -12'd193,  12'd138,  12'd77,  12'd375,  -12'd445,  -12'd64,  12'd197,  12'd243,  12'd104,  12'd417,  12'd332,  -12'd223,  
-12'd247,  12'd55,  -12'd298,  12'd500,  -12'd294,  -12'd0,  -12'd269,  -12'd11,  12'd41,  12'd61,  -12'd354,  -12'd203,  12'd8,  -12'd138,  12'd175,  -12'd245,  
12'd364,  -12'd13,  12'd321,  -12'd32,  12'd21,  12'd78,  12'd138,  -12'd134,  12'd187,  12'd241,  12'd8,  12'd367,  12'd125,  -12'd257,  -12'd87,  12'd168,  
12'd11,  -12'd388,  12'd430,  -12'd250,  -12'd390,  -12'd331,  -12'd356,  -12'd151,  -12'd296,  12'd409,  -12'd620,  12'd469,  -12'd34,  12'd335,  12'd162,  -12'd199,  
12'd47,  12'd328,  12'd392,  -12'd230,  -12'd146,  12'd8,  -12'd286,  12'd398,  12'd271,  12'd192,  -12'd346,  12'd188,  12'd61,  12'd70,  12'd101,  12'd72,  
12'd133,  12'd172,  12'd11,  12'd458,  12'd148,  12'd593,  -12'd181,  12'd515,  12'd270,  -12'd483,  -12'd175,  -12'd515,  12'd280,  -12'd258,  12'd24,  12'd84,  
-12'd219,  -12'd240,  12'd178,  -12'd228,  12'd181,  -12'd145,  -12'd295,  -12'd39,  -12'd378,  12'd189,  12'd327,  -12'd488,  -12'd78,  -12'd254,  12'd121,  12'd149,  
-12'd69,  -12'd415,  -12'd279,  12'd302,  12'd465,  -12'd272,  -12'd167,  12'd336,  12'd80,  12'd628,  12'd360,  12'd207,  -12'd109,  12'd14,  12'd117,  12'd440,  

12'd88,  12'd146,  12'd82,  12'd118,  12'd16,  12'd41,  -12'd379,  12'd18,  12'd49,  -12'd317,  12'd149,  -12'd43,  -12'd6,  -12'd223,  -12'd21,  12'd137,  
12'd263,  -12'd21,  -12'd135,  -12'd246,  12'd191,  12'd351,  12'd18,  -12'd51,  -12'd145,  -12'd121,  -12'd273,  12'd156,  12'd336,  -12'd119,  12'd168,  12'd156,  
12'd99,  -12'd82,  12'd28,  12'd167,  12'd47,  12'd218,  -12'd41,  -12'd244,  12'd160,  12'd265,  -12'd394,  -12'd292,  -12'd219,  12'd195,  12'd124,  12'd133,  
-12'd291,  -12'd68,  -12'd289,  -12'd90,  -12'd141,  -12'd60,  -12'd98,  -12'd50,  12'd386,  12'd232,  -12'd57,  -12'd20,  -12'd16,  12'd504,  12'd335,  -12'd1,  
-12'd349,  -12'd172,  -12'd124,  12'd83,  12'd98,  -12'd6,  -12'd344,  12'd143,  12'd284,  12'd219,  12'd174,  12'd78,  -12'd295,  12'd94,  12'd178,  -12'd111,  
12'd93,  12'd27,  -12'd513,  12'd104,  -12'd161,  -12'd157,  -12'd170,  -12'd388,  12'd207,  12'd405,  12'd152,  12'd55,  12'd218,  -12'd367,  -12'd175,  -12'd64,  
-12'd18,  -12'd2,  -12'd86,  -12'd266,  12'd210,  12'd70,  -12'd330,  -12'd87,  -12'd346,  12'd243,  -12'd97,  -12'd121,  -12'd10,  12'd118,  12'd43,  12'd148,  
-12'd302,  12'd567,  12'd143,  -12'd72,  12'd18,  -12'd125,  12'd115,  -12'd215,  12'd295,  12'd369,  -12'd100,  12'd434,  -12'd178,  12'd344,  -12'd211,  12'd283,  
12'd32,  -12'd261,  12'd215,  12'd144,  -12'd65,  12'd32,  -12'd264,  -12'd73,  -12'd210,  -12'd406,  -12'd371,  12'd158,  -12'd8,  12'd275,  12'd114,  12'd242,  
-12'd145,  12'd214,  12'd332,  -12'd335,  -12'd31,  12'd220,  12'd231,  -12'd152,  12'd39,  12'd72,  12'd79,  12'd282,  -12'd62,  12'd115,  -12'd160,  -12'd153,  
-12'd242,  12'd4,  12'd99,  -12'd117,  -12'd289,  -12'd2,  12'd35,  -12'd441,  12'd133,  -12'd154,  12'd176,  12'd4,  -12'd514,  -12'd414,  -12'd340,  12'd207,  
12'd311,  12'd239,  -12'd166,  12'd52,  -12'd122,  12'd402,  12'd250,  -12'd27,  12'd478,  -12'd40,  -12'd348,  12'd5,  -12'd109,  12'd106,  -12'd321,  -12'd180,  
12'd136,  12'd287,  -12'd264,  -12'd123,  12'd278,  -12'd36,  -12'd215,  12'd100,  12'd11,  -12'd108,  -12'd344,  12'd422,  12'd349,  -12'd64,  12'd30,  -12'd301,  
-12'd127,  12'd13,  12'd186,  12'd167,  -12'd59,  -12'd236,  12'd237,  -12'd329,  12'd123,  12'd82,  -12'd24,  -12'd31,  12'd1,  12'd115,  -12'd67,  12'd111,  
12'd169,  12'd23,  -12'd353,  12'd178,  12'd319,  12'd82,  -12'd115,  -12'd250,  -12'd195,  12'd29,  -12'd347,  12'd273,  12'd187,  -12'd376,  -12'd193,  -12'd64,  
12'd209,  -12'd354,  12'd228,  12'd216,  -12'd152,  -12'd26,  12'd359,  12'd28,  12'd241,  12'd7,  12'd255,  12'd40,  -12'd165,  12'd150,  12'd11,  12'd33,  
12'd64,  -12'd248,  -12'd61,  12'd191,  12'd78,  12'd361,  12'd277,  12'd200,  12'd43,  12'd55,  12'd169,  12'd212,  -12'd115,  12'd143,  12'd209,  12'd16,  
12'd260,  12'd21,  -12'd229,  12'd350,  -12'd47,  12'd66,  12'd55,  -12'd30,  -12'd375,  12'd266,  12'd26,  12'd10,  12'd185,  -12'd279,  12'd259,  -12'd149,  
-12'd79,  -12'd354,  -12'd274,  12'd77,  12'd214,  12'd65,  12'd78,  12'd113,  -12'd24,  -12'd121,  12'd255,  12'd241,  -12'd171,  -12'd331,  12'd394,  -12'd146,  
-12'd54,  12'd19,  -12'd273,  12'd62,  12'd99,  12'd239,  -12'd71,  12'd10,  -12'd171,  12'd262,  12'd370,  12'd211,  -12'd98,  -12'd165,  12'd364,  12'd381,  
12'd72,  -12'd187,  12'd91,  12'd147,  -12'd161,  -12'd372,  -12'd228,  12'd112,  -12'd337,  12'd128,  -12'd28,  -12'd99,  -12'd222,  12'd220,  12'd234,  -12'd285,  
-12'd192,  -12'd46,  -12'd164,  -12'd278,  12'd13,  -12'd206,  -12'd239,  12'd28,  -12'd298,  -12'd64,  12'd347,  -12'd147,  12'd140,  12'd451,  12'd98,  12'd202,  
12'd40,  -12'd411,  -12'd31,  12'd443,  12'd240,  12'd328,  -12'd188,  12'd224,  -12'd483,  -12'd78,  12'd123,  12'd70,  12'd310,  -12'd154,  12'd202,  12'd205,  
-12'd261,  12'd6,  -12'd38,  12'd128,  12'd377,  -12'd37,  12'd140,  12'd165,  12'd188,  12'd358,  12'd3,  12'd324,  12'd151,  -12'd90,  -12'd112,  -12'd39,  
12'd81,  12'd584,  -12'd304,  12'd375,  12'd334,  12'd349,  12'd54,  -12'd12,  12'd394,  12'd450,  12'd138,  12'd63,  12'd49,  -12'd163,  12'd141,  12'd382,  

12'd68,  12'd145,  -12'd371,  -12'd76,  12'd56,  -12'd348,  -12'd257,  -12'd213,  12'd45,  -12'd17,  12'd64,  12'd222,  -12'd541,  -12'd453,  -12'd281,  12'd1,  
12'd305,  -12'd244,  -12'd231,  12'd463,  -12'd75,  12'd47,  -12'd456,  12'd52,  -12'd108,  12'd114,  12'd243,  -12'd219,  12'd418,  -12'd171,  12'd4,  12'd332,  
-12'd157,  12'd128,  -12'd120,  12'd131,  -12'd6,  12'd368,  -12'd285,  12'd113,  12'd382,  12'd252,  -12'd340,  12'd198,  12'd279,  -12'd848,  -12'd315,  12'd139,  
-12'd57,  -12'd29,  12'd36,  12'd58,  12'd253,  12'd51,  -12'd405,  12'd25,  -12'd274,  12'd316,  -12'd24,  12'd289,  12'd214,  -12'd364,  -12'd17,  -12'd314,  
-12'd516,  -12'd235,  12'd419,  12'd105,  12'd279,  12'd15,  -12'd31,  12'd126,  -12'd206,  12'd219,  -12'd87,  -12'd70,  -12'd278,  -12'd19,  -12'd311,  -12'd369,  
12'd14,  -12'd233,  12'd159,  12'd339,  -12'd174,  12'd438,  12'd251,  12'd8,  12'd577,  12'd219,  12'd87,  12'd156,  12'd190,  12'd6,  -12'd231,  -12'd170,  
-12'd152,  12'd659,  -12'd168,  12'd13,  -12'd51,  -12'd262,  -12'd31,  12'd241,  12'd170,  -12'd11,  -12'd138,  12'd161,  12'd181,  -12'd74,  -12'd215,  12'd307,  
-12'd419,  12'd159,  12'd47,  -12'd251,  -12'd71,  12'd257,  -12'd69,  -12'd220,  -12'd211,  -12'd181,  12'd184,  12'd270,  12'd189,  -12'd112,  -12'd292,  12'd625,  
12'd122,  12'd260,  12'd52,  -12'd233,  12'd120,  -12'd43,  12'd56,  -12'd122,  12'd334,  -12'd205,  12'd246,  12'd347,  -12'd138,  12'd319,  12'd197,  -12'd38,  
-12'd319,  -12'd172,  -12'd80,  12'd205,  -12'd40,  -12'd152,  12'd116,  -12'd157,  -12'd177,  -12'd316,  12'd15,  -12'd211,  -12'd185,  12'd9,  -12'd118,  12'd134,  
12'd338,  -12'd54,  12'd373,  12'd85,  12'd626,  -12'd5,  12'd36,  12'd149,  12'd265,  12'd94,  -12'd52,  12'd104,  -12'd79,  -12'd121,  12'd146,  12'd209,  
-12'd40,  12'd222,  -12'd148,  -12'd115,  12'd189,  -12'd24,  12'd144,  12'd187,  -12'd514,  -12'd145,  12'd344,  12'd117,  12'd20,  -12'd321,  12'd170,  -12'd316,  
12'd486,  -12'd103,  12'd450,  12'd140,  -12'd189,  -12'd100,  12'd124,  12'd66,  -12'd154,  12'd9,  12'd94,  -12'd174,  -12'd300,  12'd2,  12'd105,  -12'd347,  
12'd372,  12'd153,  12'd177,  -12'd330,  -12'd119,  -12'd96,  12'd381,  -12'd434,  12'd170,  -12'd353,  -12'd41,  12'd6,  -12'd31,  -12'd11,  -12'd259,  -12'd201,  
12'd616,  12'd245,  12'd35,  -12'd152,  -12'd41,  12'd458,  12'd223,  -12'd57,  12'd145,  -12'd180,  12'd37,  12'd134,  -12'd136,  12'd449,  -12'd181,  12'd196,  
12'd46,  12'd197,  -12'd13,  12'd181,  12'd182,  -12'd312,  -12'd175,  12'd93,  -12'd213,  -12'd81,  12'd173,  12'd371,  12'd146,  12'd152,  12'd254,  -12'd305,  
-12'd45,  12'd452,  -12'd209,  -12'd227,  12'd226,  -12'd34,  -12'd156,  12'd232,  -12'd98,  -12'd0,  -12'd100,  12'd50,  -12'd281,  -12'd429,  12'd63,  12'd317,  
-12'd3,  12'd71,  -12'd310,  -12'd13,  12'd59,  -12'd209,  -12'd168,  12'd55,  12'd409,  12'd295,  -12'd309,  12'd239,  12'd71,  12'd212,  -12'd140,  12'd111,  
12'd341,  12'd127,  12'd3,  -12'd140,  -12'd78,  -12'd376,  12'd30,  -12'd166,  12'd338,  12'd215,  12'd162,  -12'd229,  -12'd204,  12'd1,  12'd56,  -12'd99,  
-12'd271,  -12'd359,  -12'd187,  -12'd58,  -12'd14,  -12'd576,  12'd247,  -12'd112,  12'd322,  12'd99,  12'd251,  -12'd260,  12'd238,  12'd166,  -12'd254,  12'd166,  
12'd39,  -12'd37,  -12'd130,  -12'd114,  -12'd339,  -12'd44,  -12'd401,  -12'd337,  -12'd200,  12'd161,  12'd322,  -12'd97,  12'd84,  12'd346,  -12'd9,  -12'd26,  
12'd39,  -12'd20,  12'd172,  12'd51,  12'd326,  12'd47,  12'd94,  12'd13,  12'd133,  12'd132,  -12'd75,  12'd260,  -12'd103,  -12'd182,  12'd145,  12'd165,  
12'd153,  12'd46,  12'd271,  -12'd61,  -12'd14,  -12'd9,  12'd120,  12'd280,  12'd14,  -12'd287,  -12'd386,  -12'd311,  -12'd330,  -12'd17,  12'd22,  -12'd244,  
-12'd173,  -12'd122,  -12'd295,  -12'd195,  -12'd107,  12'd214,  -12'd23,  -12'd236,  12'd205,  -12'd167,  -12'd190,  12'd308,  12'd94,  12'd257,  12'd289,  -12'd207,  
-12'd107,  -12'd271,  12'd127,  12'd145,  -12'd120,  12'd63,  12'd34,  -12'd65,  -12'd379,  12'd451,  12'd96,  -12'd277,  12'd142,  12'd81,  12'd170,  -12'd36,  

-12'd61,  12'd221,  -12'd32,  12'd58,  -12'd321,  -12'd4,  12'd160,  -12'd24,  -12'd351,  -12'd54,  12'd546,  12'd372,  12'd76,  12'd50,  12'd21,  12'd200,  
-12'd385,  12'd317,  -12'd168,  12'd20,  -12'd177,  -12'd1,  12'd120,  12'd14,  -12'd27,  12'd221,  12'd230,  12'd61,  -12'd95,  -12'd490,  12'd217,  -12'd5,  
-12'd10,  12'd232,  -12'd219,  -12'd308,  12'd490,  -12'd99,  12'd83,  12'd208,  12'd139,  12'd169,  12'd224,  -12'd74,  12'd67,  -12'd722,  -12'd139,  -12'd79,  
-12'd242,  -12'd441,  12'd75,  12'd245,  -12'd29,  -12'd220,  -12'd166,  12'd293,  12'd26,  -12'd64,  -12'd41,  12'd254,  -12'd321,  12'd78,  -12'd128,  -12'd68,  
-12'd117,  -12'd320,  12'd251,  -12'd75,  -12'd315,  -12'd261,  -12'd48,  -12'd30,  -12'd19,  12'd67,  -12'd124,  12'd25,  -12'd11,  -12'd133,  -12'd87,  12'd292,  
12'd107,  12'd398,  -12'd190,  12'd37,  -12'd94,  12'd100,  -12'd352,  -12'd98,  -12'd31,  -12'd379,  12'd188,  -12'd3,  12'd338,  12'd267,  12'd213,  12'd424,  
12'd312,  12'd46,  -12'd191,  -12'd289,  12'd133,  -12'd34,  12'd182,  -12'd144,  12'd297,  -12'd372,  12'd137,  12'd214,  12'd27,  -12'd50,  12'd323,  12'd99,  
12'd280,  12'd212,  -12'd324,  12'd36,  12'd287,  -12'd114,  12'd98,  12'd277,  12'd249,  12'd112,  -12'd178,  12'd578,  -12'd303,  -12'd85,  -12'd126,  12'd285,  
12'd112,  12'd119,  -12'd396,  -12'd67,  12'd143,  12'd53,  12'd430,  -12'd117,  -12'd37,  -12'd9,  -12'd257,  -12'd13,  12'd36,  -12'd96,  12'd58,  12'd88,  
-12'd384,  -12'd386,  -12'd209,  12'd113,  12'd89,  -12'd102,  12'd322,  -12'd9,  12'd114,  -12'd63,  -12'd20,  -12'd76,  12'd37,  12'd217,  -12'd328,  12'd47,  
-12'd168,  -12'd160,  12'd304,  12'd139,  -12'd100,  -12'd30,  12'd303,  -12'd204,  -12'd207,  -12'd88,  -12'd129,  -12'd250,  -12'd28,  -12'd24,  -12'd166,  -12'd291,  
12'd270,  -12'd69,  -12'd253,  12'd58,  -12'd55,  -12'd301,  -12'd295,  -12'd201,  -12'd291,  -12'd280,  -12'd13,  -12'd145,  12'd38,  12'd254,  12'd359,  12'd24,  
12'd180,  12'd1,  12'd176,  12'd47,  12'd123,  -12'd250,  -12'd58,  -12'd296,  -12'd104,  12'd17,  12'd246,  12'd82,  -12'd79,  12'd20,  -12'd141,  -12'd23,  
12'd260,  -12'd406,  -12'd110,  -12'd313,  12'd157,  12'd176,  -12'd304,  -12'd23,  12'd30,  -12'd10,  12'd146,  -12'd4,  -12'd63,  -12'd41,  12'd110,  12'd71,  
-12'd389,  -12'd33,  12'd183,  12'd109,  12'd231,  12'd241,  12'd3,  -12'd214,  -12'd2,  12'd342,  -12'd86,  12'd225,  -12'd173,  12'd7,  -12'd269,  -12'd11,  
12'd205,  12'd310,  12'd245,  12'd136,  12'd21,  -12'd11,  -12'd109,  -12'd148,  12'd324,  12'd218,  -12'd133,  -12'd585,  12'd88,  -12'd118,  -12'd272,  -12'd108,  
-12'd253,  12'd36,  -12'd346,  -12'd128,  12'd307,  -12'd153,  12'd130,  12'd21,  -12'd70,  -12'd9,  12'd64,  -12'd94,  12'd105,  -12'd112,  -12'd389,  -12'd317,  
12'd47,  -12'd52,  12'd95,  -12'd149,  -12'd275,  -12'd262,  12'd48,  12'd375,  12'd56,  12'd20,  -12'd19,  -12'd258,  12'd206,  12'd274,  -12'd135,  12'd249,  
12'd339,  -12'd89,  12'd208,  12'd239,  12'd32,  12'd40,  -12'd338,  -12'd244,  -12'd164,  12'd97,  12'd216,  12'd300,  -12'd244,  12'd348,  12'd278,  12'd144,  
12'd252,  12'd356,  -12'd428,  12'd206,  -12'd101,  12'd120,  12'd163,  12'd331,  -12'd74,  12'd318,  -12'd48,  -12'd245,  12'd187,  12'd23,  12'd127,  -12'd159,  
12'd185,  12'd85,  -12'd223,  12'd28,  -12'd109,  -12'd245,  12'd124,  -12'd335,  12'd243,  -12'd78,  12'd210,  12'd0,  12'd20,  -12'd496,  12'd180,  12'd192,  
12'd280,  12'd327,  12'd66,  -12'd272,  -12'd442,  -12'd196,  12'd196,  -12'd460,  12'd568,  -12'd231,  -12'd357,  -12'd86,  -12'd165,  -12'd292,  -12'd338,  12'd173,  
-12'd287,  12'd114,  12'd260,  -12'd210,  -12'd129,  12'd119,  12'd7,  -12'd76,  12'd522,  12'd702,  -12'd370,  12'd149,  12'd7,  12'd651,  12'd219,  -12'd40,  
12'd256,  -12'd251,  12'd93,  -12'd26,  -12'd85,  12'd10,  12'd196,  12'd280,  12'd354,  -12'd200,  -12'd242,  12'd349,  -12'd12,  12'd396,  -12'd291,  -12'd164,  
-12'd196,  12'd330,  12'd449,  12'd354,  12'd95,  -12'd101,  12'd414,  12'd351,  12'd349,  -12'd90,  -12'd339,  -12'd27,  12'd206,  12'd85,  12'd93,  12'd33,  

-12'd206,  -12'd144,  -12'd209,  12'd162,  12'd243,  -12'd154,  -12'd723,  12'd111,  -12'd190,  -12'd65,  -12'd269,  -12'd31,  12'd165,  -12'd97,  12'd360,  12'd271,  
-12'd179,  -12'd90,  -12'd82,  12'd85,  -12'd146,  -12'd237,  -12'd22,  12'd398,  -12'd83,  12'd369,  -12'd114,  -12'd78,  12'd77,  -12'd424,  -12'd128,  -12'd23,  
-12'd212,  12'd242,  12'd138,  12'd484,  12'd27,  -12'd235,  -12'd317,  12'd381,  -12'd251,  -12'd165,  -12'd360,  12'd105,  12'd99,  -12'd616,  -12'd41,  12'd363,  
12'd125,  -12'd152,  -12'd159,  12'd236,  -12'd116,  12'd248,  -12'd137,  12'd134,  -12'd15,  12'd210,  12'd250,  12'd83,  12'd290,  -12'd300,  -12'd44,  12'd571,  
-12'd84,  -12'd435,  12'd83,  12'd24,  12'd12,  12'd42,  12'd300,  -12'd218,  12'd209,  12'd535,  12'd83,  12'd170,  12'd174,  -12'd122,  -12'd99,  12'd49,  
-12'd260,  12'd151,  12'd24,  12'd251,  12'd279,  12'd29,  -12'd349,  -12'd250,  12'd162,  12'd116,  -12'd204,  12'd384,  12'd336,  -12'd374,  -12'd460,  12'd241,  
-12'd147,  -12'd34,  -12'd124,  -12'd88,  12'd131,  12'd21,  12'd157,  -12'd20,  -12'd13,  -12'd235,  12'd96,  -12'd199,  12'd217,  -12'd363,  -12'd338,  12'd103,  
-12'd6,  12'd63,  -12'd199,  12'd170,  12'd71,  -12'd37,  12'd140,  -12'd90,  -12'd413,  12'd364,  12'd177,  -12'd189,  12'd177,  12'd521,  12'd25,  12'd205,  
12'd51,  12'd84,  12'd527,  -12'd212,  -12'd30,  12'd261,  12'd103,  -12'd90,  -12'd186,  12'd71,  12'd72,  12'd270,  12'd29,  12'd174,  12'd240,  12'd577,  
12'd1,  -12'd39,  -12'd255,  12'd192,  12'd6,  12'd169,  12'd343,  12'd195,  12'd27,  -12'd101,  -12'd103,  12'd11,  -12'd14,  12'd208,  12'd66,  -12'd116,  
-12'd272,  12'd271,  -12'd327,  12'd107,  -12'd74,  -12'd55,  12'd31,  12'd210,  12'd428,  -12'd392,  12'd70,  12'd32,  -12'd150,  -12'd362,  -12'd246,  12'd138,  
12'd78,  -12'd365,  -12'd167,  -12'd516,  12'd384,  12'd0,  12'd65,  -12'd70,  12'd47,  -12'd114,  -12'd6,  -12'd157,  12'd302,  -12'd65,  12'd130,  12'd69,  
-12'd138,  -12'd182,  12'd345,  12'd162,  12'd193,  12'd9,  -12'd159,  -12'd383,  -12'd182,  -12'd64,  -12'd301,  12'd11,  -12'd209,  12'd196,  12'd196,  -12'd154,  
12'd203,  12'd318,  12'd122,  -12'd157,  12'd407,  12'd343,  12'd183,  12'd364,  12'd233,  12'd291,  12'd55,  12'd179,  12'd323,  12'd105,  -12'd69,  12'd5,  
12'd423,  -12'd102,  12'd374,  -12'd1,  12'd205,  12'd276,  12'd260,  12'd76,  -12'd313,  -12'd295,  -12'd63,  12'd271,  12'd234,  12'd15,  12'd224,  12'd138,  
12'd89,  12'd37,  -12'd40,  12'd215,  -12'd224,  -12'd119,  12'd107,  12'd179,  12'd146,  12'd88,  -12'd196,  12'd138,  -12'd301,  -12'd120,  12'd114,  12'd54,  
12'd357,  12'd10,  -12'd9,  -12'd148,  -12'd92,  12'd159,  -12'd244,  12'd3,  12'd196,  12'd103,  12'd68,  -12'd100,  12'd4,  12'd153,  -12'd1,  -12'd185,  
-12'd173,  12'd61,  12'd151,  12'd278,  12'd19,  -12'd271,  12'd36,  12'd289,  12'd35,  -12'd348,  12'd287,  -12'd96,  -12'd56,  -12'd84,  -12'd8,  -12'd109,  
-12'd368,  -12'd314,  12'd31,  12'd24,  -12'd144,  -12'd169,  12'd261,  -12'd129,  -12'd252,  -12'd277,  12'd394,  12'd241,  12'd208,  12'd10,  12'd317,  -12'd68,  
12'd159,  -12'd40,  -12'd70,  -12'd393,  12'd132,  12'd63,  12'd201,  -12'd162,  -12'd339,  -12'd97,  12'd290,  -12'd24,  -12'd35,  -12'd266,  -12'd119,  12'd162,  
-12'd86,  12'd38,  -12'd8,  -12'd89,  12'd3,  -12'd185,  -12'd118,  -12'd17,  -12'd314,  12'd7,  -12'd31,  -12'd37,  -12'd223,  -12'd234,  12'd335,  12'd107,  
-12'd87,  12'd123,  -12'd131,  -12'd61,  -12'd68,  -12'd360,  -12'd9,  -12'd393,  12'd150,  -12'd342,  -12'd54,  12'd97,  12'd192,  12'd95,  -12'd281,  12'd243,  
12'd31,  12'd124,  12'd118,  -12'd378,  -12'd339,  -12'd394,  -12'd46,  12'd200,  -12'd21,  12'd419,  -12'd407,  12'd186,  -12'd270,  12'd105,  -12'd331,  -12'd13,  
-12'd165,  12'd155,  12'd202,  -12'd164,  12'd161,  -12'd50,  12'd215,  -12'd127,  -12'd312,  -12'd57,  12'd17,  12'd100,  -12'd291,  -12'd302,  12'd121,  -12'd257,  
12'd103,  12'd206,  12'd3,  -12'd398,  12'd7,  -12'd443,  -12'd141,  -12'd56,  -12'd300,  -12'd171,  12'd136,  -12'd567,  -12'd228,  -12'd156,  -12'd438,  -12'd89,  

-12'd207,  12'd291,  -12'd54,  12'd77,  12'd206,  12'd213,  -12'd197,  -12'd22,  12'd377,  12'd82,  12'd65,  -12'd288,  -12'd72,  12'd156,  -12'd124,  -12'd191,  
-12'd264,  -12'd105,  12'd446,  12'd331,  12'd144,  12'd117,  12'd146,  12'd21,  -12'd98,  -12'd100,  -12'd166,  12'd4,  12'd394,  12'd98,  12'd379,  12'd379,  
12'd189,  -12'd317,  12'd229,  -12'd205,  -12'd28,  12'd120,  12'd378,  12'd107,  12'd123,  12'd321,  12'd237,  12'd224,  -12'd91,  12'd353,  12'd274,  -12'd195,  
12'd199,  -12'd113,  -12'd75,  12'd308,  -12'd181,  -12'd51,  12'd135,  -12'd280,  12'd444,  12'd45,  12'd128,  -12'd226,  -12'd83,  12'd394,  -12'd520,  -12'd139,  
12'd107,  -12'd82,  -12'd286,  -12'd384,  12'd264,  -12'd287,  12'd373,  12'd67,  12'd15,  -12'd167,  12'd248,  -12'd102,  12'd144,  -12'd177,  -12'd250,  -12'd142,  
-12'd364,  -12'd197,  -12'd117,  -12'd427,  12'd341,  -12'd269,  12'd101,  12'd208,  -12'd214,  12'd90,  12'd75,  -12'd426,  -12'd233,  -12'd304,  12'd37,  12'd29,  
-12'd188,  -12'd179,  12'd39,  12'd127,  -12'd76,  -12'd220,  -12'd682,  -12'd128,  -12'd317,  12'd302,  -12'd153,  -12'd325,  -12'd173,  -12'd547,  12'd11,  12'd8,  
12'd227,  -12'd647,  12'd398,  12'd124,  -12'd21,  12'd355,  12'd32,  12'd8,  -12'd777,  12'd21,  12'd45,  -12'd91,  -12'd157,  12'd91,  12'd196,  12'd88,  
12'd432,  -12'd200,  12'd349,  12'd203,  12'd42,  -12'd166,  12'd273,  12'd534,  -12'd436,  -12'd72,  12'd239,  -12'd289,  -12'd151,  12'd288,  12'd34,  -12'd29,  
12'd610,  -12'd262,  12'd216,  12'd269,  -12'd151,  -12'd31,  -12'd171,  -12'd80,  12'd203,  12'd229,  12'd145,  -12'd316,  -12'd67,  12'd100,  -12'd339,  -12'd7,  
-12'd363,  -12'd129,  -12'd506,  -12'd2,  12'd201,  -12'd293,  -12'd120,  12'd121,  12'd250,  12'd40,  -12'd74,  -12'd617,  12'd73,  -12'd649,  -12'd165,  -12'd295,  
-12'd23,  -12'd176,  -12'd139,  12'd122,  -12'd405,  12'd34,  -12'd405,  -12'd127,  12'd74,  12'd85,  12'd51,  12'd75,  -12'd404,  -12'd36,  12'd190,  12'd165,  
12'd458,  12'd195,  12'd317,  12'd56,  -12'd434,  12'd8,  -12'd392,  12'd128,  -12'd128,  12'd416,  12'd250,  -12'd115,  12'd130,  -12'd53,  12'd508,  12'd190,  
12'd174,  -12'd222,  12'd78,  12'd66,  -12'd57,  12'd43,  -12'd170,  12'd222,  -12'd271,  12'd272,  -12'd141,  -12'd324,  12'd499,  -12'd258,  -12'd209,  12'd122,  
-12'd256,  -12'd190,  -12'd24,  12'd192,  -12'd295,  -12'd281,  12'd161,  12'd129,  12'd271,  -12'd65,  12'd218,  -12'd49,  -12'd62,  12'd40,  -12'd157,  -12'd8,  
-12'd509,  -12'd22,  -12'd253,  12'd89,  12'd49,  12'd102,  12'd27,  12'd143,  12'd133,  12'd230,  12'd156,  -12'd446,  -12'd331,  12'd194,  12'd66,  -12'd163,  
12'd185,  12'd249,  -12'd126,  -12'd54,  -12'd234,  12'd306,  12'd98,  -12'd24,  -12'd264,  12'd115,  12'd72,  -12'd44,  12'd113,  -12'd55,  12'd108,  -12'd148,  
12'd153,  -12'd7,  -12'd297,  12'd177,  -12'd139,  -12'd17,  12'd124,  12'd183,  -12'd42,  12'd87,  12'd161,  12'd56,  12'd306,  -12'd376,  12'd108,  12'd169,  
-12'd3,  -12'd149,  12'd379,  12'd101,  -12'd245,  -12'd154,  -12'd229,  -12'd93,  -12'd183,  12'd57,  12'd231,  12'd32,  -12'd188,  -12'd53,  12'd7,  12'd10,  
-12'd204,  -12'd67,  12'd2,  -12'd59,  12'd75,  -12'd104,  12'd60,  12'd272,  -12'd186,  12'd318,  -12'd31,  -12'd100,  -12'd24,  12'd170,  -12'd191,  -12'd62,  
12'd106,  12'd369,  -12'd111,  12'd220,  -12'd51,  12'd191,  12'd259,  -12'd112,  12'd233,  -12'd64,  -12'd175,  12'd316,  12'd83,  -12'd137,  12'd109,  -12'd42,  
12'd14,  12'd265,  12'd85,  -12'd31,  12'd85,  -12'd21,  12'd126,  12'd102,  -12'd148,  -12'd68,  -12'd273,  12'd27,  12'd86,  12'd237,  12'd251,  -12'd163,  
12'd178,  -12'd104,  12'd122,  -12'd169,  12'd178,  12'd147,  12'd131,  -12'd138,  12'd175,  12'd275,  12'd190,  -12'd40,  -12'd162,  -12'd222,  12'd208,  12'd180,  
-12'd117,  12'd135,  -12'd20,  -12'd188,  -12'd238,  -12'd403,  12'd263,  -12'd255,  -12'd237,  -12'd168,  12'd71,  12'd60,  -12'd225,  12'd440,  12'd132,  12'd138,  
12'd159,  12'd353,  -12'd20,  12'd177,  12'd128,  -12'd334,  -12'd219,  -12'd147,  12'd369,  -12'd208,  12'd132,  -12'd63,  -12'd456,  12'd320,  -12'd226,  -12'd23,  

-12'd334,  12'd207,  -12'd142,  -12'd203,  -12'd98,  12'd0,  -12'd86,  -12'd329,  -12'd231,  -12'd351,  -12'd532,  -12'd249,  -12'd170,  -12'd324,  -12'd217,  -12'd219,  
-12'd280,  12'd233,  -12'd63,  12'd274,  -12'd67,  12'd410,  12'd95,  12'd86,  12'd178,  -12'd65,  -12'd591,  12'd68,  -12'd263,  12'd126,  12'd29,  12'd101,  
12'd233,  -12'd33,  -12'd127,  12'd43,  12'd456,  12'd322,  12'd248,  -12'd288,  -12'd389,  -12'd239,  12'd232,  12'd173,  -12'd279,  -12'd182,  12'd187,  -12'd370,  
-12'd227,  -12'd97,  -12'd19,  12'd301,  -12'd24,  12'd309,  -12'd191,  -12'd57,  -12'd85,  -12'd114,  12'd171,  -12'd157,  12'd384,  12'd631,  -12'd164,  -12'd334,  
-12'd229,  -12'd367,  -12'd109,  12'd289,  12'd361,  -12'd79,  12'd112,  12'd20,  -12'd351,  12'd181,  -12'd152,  -12'd343,  -12'd194,  -12'd99,  12'd151,  -12'd393,  
-12'd231,  -12'd138,  -12'd415,  12'd75,  12'd431,  -12'd427,  -12'd88,  -12'd404,  12'd80,  -12'd122,  -12'd33,  12'd171,  -12'd94,  -12'd30,  -12'd373,  -12'd438,  
12'd203,  -12'd54,  12'd175,  -12'd404,  12'd275,  -12'd152,  -12'd104,  -12'd178,  -12'd241,  12'd110,  -12'd286,  -12'd447,  -12'd481,  -12'd252,  -12'd103,  -12'd397,  
12'd173,  12'd314,  12'd212,  12'd10,  -12'd468,  12'd36,  -12'd44,  12'd123,  12'd231,  12'd168,  -12'd94,  -12'd193,  -12'd147,  12'd157,  12'd232,  -12'd310,  
12'd13,  12'd6,  12'd279,  12'd73,  -12'd51,  -12'd179,  12'd318,  -12'd144,  -12'd157,  -12'd147,  12'd223,  12'd302,  12'd98,  12'd617,  12'd188,  12'd184,  
-12'd174,  12'd127,  12'd150,  -12'd138,  -12'd8,  -12'd93,  12'd155,  -12'd289,  12'd92,  -12'd85,  -12'd22,  12'd60,  -12'd143,  -12'd61,  -12'd326,  -12'd257,  
-12'd343,  -12'd296,  -12'd8,  12'd160,  12'd38,  -12'd160,  -12'd34,  12'd57,  12'd351,  -12'd147,  12'd124,  -12'd110,  -12'd71,  12'd156,  -12'd35,  -12'd331,  
-12'd84,  -12'd277,  12'd24,  12'd225,  12'd172,  12'd381,  12'd80,  -12'd66,  12'd223,  -12'd66,  -12'd74,  -12'd202,  12'd59,  -12'd157,  12'd91,  12'd115,  
12'd229,  12'd27,  12'd201,  -12'd197,  12'd163,  12'd404,  -12'd20,  12'd281,  12'd297,  -12'd58,  -12'd293,  12'd224,  -12'd0,  12'd62,  12'd207,  -12'd320,  
12'd144,  -12'd125,  12'd121,  -12'd44,  -12'd6,  12'd132,  12'd163,  12'd140,  12'd289,  12'd52,  -12'd182,  -12'd23,  12'd240,  12'd260,  12'd144,  -12'd195,  
12'd209,  12'd318,  -12'd33,  12'd119,  12'd55,  -12'd476,  -12'd194,  -12'd8,  -12'd356,  -12'd497,  12'd67,  -12'd228,  -12'd132,  -12'd202,  -12'd8,  12'd31,  
12'd198,  -12'd95,  12'd208,  12'd64,  -12'd148,  -12'd245,  12'd285,  -12'd280,  12'd78,  -12'd492,  12'd567,  12'd314,  12'd118,  -12'd126,  -12'd84,  12'd162,  
12'd112,  -12'd96,  -12'd3,  -12'd236,  -12'd608,  12'd56,  12'd278,  -12'd26,  12'd102,  12'd88,  12'd267,  -12'd297,  12'd209,  12'd309,  12'd98,  12'd398,  
12'd196,  -12'd202,  -12'd215,  12'd239,  -12'd211,  12'd292,  12'd69,  12'd454,  12'd277,  -12'd195,  12'd284,  -12'd227,  12'd121,  12'd300,  12'd324,  12'd96,  
-12'd85,  -12'd188,  -12'd234,  -12'd12,  -12'd91,  12'd58,  12'd177,  12'd347,  -12'd185,  12'd236,  -12'd18,  12'd34,  -12'd78,  12'd344,  -12'd84,  -12'd63,  
12'd278,  12'd159,  -12'd96,  12'd81,  -12'd615,  -12'd182,  -12'd519,  -12'd315,  -12'd531,  -12'd578,  12'd108,  12'd163,  -12'd414,  12'd429,  -12'd103,  -12'd193,  
12'd67,  -12'd467,  12'd43,  -12'd273,  -12'd303,  12'd67,  12'd389,  -12'd138,  12'd69,  12'd97,  12'd127,  -12'd1,  -12'd222,  12'd236,  12'd5,  -12'd189,  
12'd225,  12'd97,  -12'd22,  -12'd337,  12'd85,  12'd117,  12'd430,  -12'd356,  12'd494,  12'd375,  12'd11,  -12'd39,  -12'd328,  12'd4,  -12'd127,  12'd86,  
12'd31,  -12'd132,  12'd539,  -12'd320,  12'd218,  -12'd152,  -12'd65,  12'd162,  12'd254,  12'd249,  -12'd305,  12'd51,  -12'd254,  12'd276,  12'd215,  -12'd250,  
-12'd576,  -12'd295,  -12'd105,  12'd196,  12'd361,  -12'd95,  12'd306,  -12'd38,  12'd22,  12'd106,  -12'd170,  -12'd307,  12'd24,  -12'd82,  12'd37,  -12'd257,  
12'd2,  12'd129,  12'd415,  12'd106,  -12'd6,  12'd92,  -12'd206,  12'd62,  12'd18,  12'd177,  -12'd313,  12'd135,  12'd393,  12'd41,  -12'd199,  12'd55,  

-12'd229,  -12'd106,  -12'd296,  12'd315,  12'd269,  -12'd182,  12'd88,  12'd203,  -12'd333,  -12'd244,  12'd370,  -12'd486,  12'd132,  -12'd309,  -12'd213,  12'd10,  
12'd56,  -12'd134,  -12'd208,  12'd300,  12'd82,  12'd208,  -12'd94,  12'd138,  12'd46,  -12'd137,  -12'd321,  -12'd17,  12'd336,  -12'd525,  -12'd139,  -12'd218,  
-12'd195,  -12'd266,  -12'd314,  12'd139,  -12'd3,  -12'd122,  -12'd395,  -12'd24,  -12'd235,  -12'd149,  12'd170,  -12'd401,  -12'd126,  -12'd324,  -12'd217,  12'd116,  
-12'd215,  -12'd532,  12'd251,  12'd258,  12'd196,  -12'd5,  12'd64,  -12'd148,  -12'd143,  12'd321,  12'd100,  -12'd47,  -12'd120,  -12'd200,  12'd332,  12'd241,  
-12'd226,  -12'd437,  12'd155,  -12'd56,  -12'd61,  -12'd45,  -12'd28,  -12'd255,  12'd277,  -12'd244,  -12'd53,  -12'd5,  -12'd385,  12'd14,  -12'd9,  -12'd59,  
-12'd215,  12'd48,  -12'd454,  12'd7,  -12'd312,  -12'd404,  12'd10,  -12'd164,  -12'd51,  -12'd117,  12'd487,  -12'd161,  12'd108,  12'd31,  -12'd206,  -12'd362,  
-12'd98,  -12'd310,  -12'd142,  12'd96,  12'd193,  -12'd384,  12'd161,  -12'd312,  -12'd88,  12'd143,  -12'd94,  12'd436,  -12'd203,  -12'd427,  12'd226,  12'd90,  
-12'd43,  12'd137,  -12'd97,  12'd41,  12'd361,  12'd149,  12'd119,  -12'd52,  12'd86,  12'd219,  12'd108,  12'd349,  12'd217,  12'd11,  12'd97,  12'd234,  
12'd254,  -12'd219,  -12'd344,  -12'd85,  12'd431,  12'd69,  -12'd13,  12'd231,  -12'd63,  12'd239,  12'd1,  12'd452,  12'd28,  12'd46,  -12'd29,  12'd49,  
-12'd286,  12'd267,  12'd291,  12'd405,  -12'd19,  12'd41,  12'd421,  12'd75,  12'd130,  12'd384,  12'd74,  12'd302,  -12'd73,  -12'd113,  12'd313,  12'd50,  
-12'd215,  12'd230,  12'd292,  12'd201,  -12'd207,  12'd41,  -12'd207,  -12'd164,  12'd62,  -12'd168,  12'd54,  -12'd121,  -12'd237,  -12'd370,  -12'd322,  -12'd248,  
12'd6,  -12'd31,  -12'd44,  -12'd150,  -12'd169,  -12'd46,  -12'd356,  12'd61,  -12'd28,  12'd103,  -12'd339,  12'd95,  -12'd254,  -12'd556,  -12'd121,  -12'd44,  
12'd399,  -12'd387,  -12'd131,  -12'd211,  -12'd123,  -12'd475,  -12'd196,  -12'd6,  12'd89,  12'd190,  12'd89,  -12'd64,  -12'd77,  -12'd210,  12'd314,  12'd238,  
-12'd156,  -12'd60,  12'd123,  -12'd220,  12'd221,  12'd125,  12'd45,  12'd259,  -12'd238,  12'd44,  12'd248,  -12'd67,  12'd119,  -12'd221,  -12'd18,  12'd153,  
-12'd39,  -12'd180,  -12'd9,  12'd270,  12'd283,  12'd22,  -12'd109,  12'd292,  12'd23,  12'd7,  -12'd84,  12'd265,  -12'd223,  12'd40,  12'd0,  -12'd17,  
-12'd211,  -12'd159,  12'd47,  -12'd20,  -12'd261,  12'd260,  -12'd511,  12'd190,  12'd294,  12'd13,  -12'd170,  -12'd274,  12'd348,  12'd259,  -12'd262,  12'd94,  
-12'd59,  -12'd478,  -12'd359,  12'd132,  -12'd11,  -12'd160,  -12'd272,  12'd333,  -12'd333,  12'd215,  12'd267,  12'd146,  12'd170,  -12'd56,  -12'd16,  12'd165,  
-12'd359,  12'd134,  -12'd138,  -12'd163,  12'd255,  -12'd324,  -12'd31,  12'd184,  -12'd187,  -12'd237,  12'd34,  -12'd190,  12'd193,  -12'd213,  12'd255,  -12'd225,  
12'd148,  12'd205,  12'd170,  12'd24,  12'd334,  12'd132,  -12'd124,  -12'd113,  -12'd105,  12'd213,  -12'd108,  12'd95,  -12'd148,  12'd51,  12'd134,  12'd152,  
12'd55,  -12'd67,  12'd238,  -12'd156,  -12'd23,  -12'd80,  12'd229,  12'd10,  -12'd177,  12'd288,  12'd237,  -12'd203,  12'd389,  -12'd107,  12'd141,  -12'd41,  
-12'd190,  -12'd17,  12'd114,  -12'd59,  12'd10,  12'd111,  -12'd284,  12'd76,  12'd71,  12'd112,  -12'd24,  -12'd101,  12'd144,  12'd56,  12'd291,  -12'd112,  
12'd2,  12'd29,  12'd27,  12'd198,  12'd226,  -12'd30,  12'd302,  -12'd261,  -12'd447,  -12'd268,  -12'd5,  12'd338,  12'd78,  -12'd289,  -12'd183,  12'd0,  
-12'd32,  12'd35,  12'd50,  12'd41,  12'd301,  12'd89,  -12'd18,  -12'd276,  -12'd45,  12'd163,  -12'd123,  12'd401,  12'd355,  -12'd223,  -12'd23,  12'd297,  
12'd239,  12'd385,  -12'd190,  -12'd173,  12'd143,  12'd99,  12'd63,  -12'd326,  12'd250,  -12'd11,  -12'd47,  -12'd197,  12'd197,  -12'd102,  -12'd181,  12'd318,  
12'd387,  12'd591,  12'd210,  -12'd42,  12'd286,  12'd251,  -12'd65,  12'd328,  12'd531,  12'd751,  -12'd154,  12'd371,  -12'd331,  12'd397,  12'd107,  12'd201,  

12'd84,  12'd72,  12'd442,  12'd84,  -12'd63,  12'd75,  12'd206,  -12'd100,  12'd158,  12'd235,  -12'd97,  -12'd89,  12'd80,  12'd134,  -12'd311,  12'd177,  
-12'd30,  -12'd80,  12'd101,  -12'd154,  -12'd196,  12'd7,  12'd126,  -12'd121,  -12'd187,  -12'd52,  12'd361,  12'd8,  -12'd168,  12'd623,  -12'd386,  12'd53,  
-12'd128,  -12'd467,  12'd281,  -12'd103,  -12'd435,  -12'd107,  12'd234,  12'd201,  -12'd94,  12'd224,  12'd306,  -12'd224,  12'd351,  12'd404,  -12'd216,  -12'd354,  
12'd343,  12'd422,  -12'd140,  12'd33,  12'd99,  -12'd136,  12'd183,  12'd179,  -12'd2,  -12'd68,  12'd279,  12'd369,  12'd22,  -12'd42,  -12'd189,  -12'd102,  
12'd700,  12'd514,  -12'd219,  12'd200,  -12'd128,  12'd392,  -12'd49,  12'd91,  -12'd267,  12'd66,  -12'd14,  12'd346,  12'd229,  12'd77,  12'd150,  12'd38,  
12'd51,  12'd21,  12'd31,  12'd147,  -12'd151,  12'd331,  12'd365,  12'd8,  12'd74,  -12'd72,  12'd32,  12'd5,  -12'd55,  12'd246,  12'd355,  -12'd105,  
12'd101,  -12'd381,  -12'd104,  12'd170,  -12'd1,  12'd165,  12'd191,  12'd137,  12'd74,  -12'd221,  12'd530,  12'd16,  -12'd153,  12'd21,  12'd216,  -12'd347,  
-12'd292,  -12'd113,  -12'd115,  -12'd87,  -12'd540,  -12'd8,  -12'd84,  -12'd340,  12'd126,  12'd18,  12'd187,  -12'd511,  12'd219,  12'd125,  -12'd127,  -12'd267,  
-12'd55,  -12'd66,  -12'd441,  12'd203,  12'd154,  -12'd343,  -12'd179,  12'd115,  -12'd7,  12'd75,  12'd140,  12'd48,  12'd145,  -12'd6,  -12'd172,  -12'd163,  
12'd90,  -12'd474,  -12'd311,  12'd125,  12'd22,  12'd288,  -12'd403,  -12'd211,  12'd150,  12'd73,  -12'd92,  12'd201,  -12'd22,  -12'd59,  -12'd263,  12'd468,  
-12'd206,  12'd152,  12'd124,  12'd228,  -12'd2,  12'd172,  12'd118,  12'd148,  -12'd253,  -12'd235,  -12'd15,  12'd72,  12'd378,  12'd209,  12'd383,  12'd89,  
12'd140,  -12'd257,  12'd65,  12'd50,  12'd336,  12'd52,  -12'd31,  12'd297,  12'd83,  -12'd167,  12'd519,  12'd123,  -12'd34,  -12'd302,  -12'd46,  12'd162,  
-12'd143,  -12'd120,  -12'd228,  12'd220,  -12'd128,  -12'd337,  12'd2,  -12'd103,  -12'd129,  12'd346,  12'd161,  -12'd76,  -12'd201,  12'd16,  -12'd471,  -12'd52,  
-12'd186,  12'd45,  -12'd227,  12'd273,  12'd433,  12'd71,  12'd70,  -12'd162,  12'd39,  12'd225,  12'd115,  12'd19,  -12'd142,  12'd203,  12'd205,  12'd3,  
-12'd372,  -12'd75,  12'd169,  12'd300,  -12'd35,  -12'd314,  -12'd338,  -12'd159,  12'd128,  12'd411,  12'd44,  -12'd258,  -12'd238,  -12'd79,  12'd110,  12'd80,  
-12'd104,  12'd191,  -12'd208,  12'd274,  12'd256,  -12'd150,  12'd72,  12'd322,  12'd26,  -12'd15,  -12'd3,  -12'd433,  12'd315,  -12'd53,  -12'd58,  12'd464,  
-12'd464,  12'd408,  -12'd80,  12'd177,  12'd159,  -12'd53,  12'd14,  -12'd1,  -12'd96,  -12'd280,  -12'd431,  12'd268,  12'd177,  -12'd373,  -12'd205,  12'd71,  
-12'd293,  -12'd145,  -12'd295,  -12'd183,  12'd253,  12'd190,  -12'd72,  -12'd74,  12'd57,  12'd200,  12'd110,  12'd361,  12'd194,  12'd405,  -12'd10,  12'd363,  
12'd45,  -12'd381,  12'd30,  -12'd137,  12'd291,  12'd1,  12'd87,  12'd45,  12'd161,  12'd43,  12'd225,  12'd362,  12'd76,  12'd31,  -12'd90,  12'd360,  
-12'd230,  12'd1,  12'd391,  -12'd138,  12'd284,  12'd22,  12'd361,  -12'd25,  12'd29,  12'd168,  12'd46,  -12'd148,  -12'd159,  12'd77,  -12'd195,  12'd64,  
12'd199,  -12'd105,  -12'd332,  -12'd360,  12'd151,  -12'd96,  12'd306,  -12'd174,  12'd181,  12'd77,  12'd76,  12'd244,  -12'd171,  -12'd483,  -12'd162,  12'd83,  
12'd112,  12'd310,  -12'd94,  -12'd309,  12'd391,  12'd115,  12'd396,  12'd159,  12'd82,  -12'd219,  -12'd228,  -12'd67,  12'd89,  -12'd138,  -12'd90,  12'd56,  
-12'd153,  12'd37,  12'd168,  -12'd86,  12'd277,  -12'd437,  12'd237,  -12'd116,  12'd205,  12'd207,  -12'd117,  12'd147,  12'd58,  12'd29,  12'd297,  12'd37,  
12'd283,  -12'd83,  12'd381,  -12'd24,  12'd18,  -12'd328,  -12'd154,  12'd46,  -12'd26,  12'd258,  12'd191,  -12'd185,  12'd190,  12'd469,  -12'd104,  -12'd47,  
12'd289,  -12'd44,  -12'd169,  -12'd80,  -12'd95,  12'd465,  12'd48,  12'd195,  -12'd49,  -12'd11,  -12'd170,  12'd126,  -12'd161,  12'd219,  12'd471,  -12'd130,  

-12'd413,  -12'd460,  -12'd162,  -12'd157,  12'd124,  -12'd113,  -12'd382,  -12'd94,  12'd78,  12'd94,  -12'd350,  -12'd200,  -12'd510,  -12'd379,  12'd129,  -12'd56,  
12'd179,  -12'd88,  12'd162,  -12'd130,  -12'd61,  12'd288,  12'd30,  -12'd52,  -12'd205,  -12'd49,  -12'd328,  12'd371,  12'd206,  12'd270,  -12'd250,  -12'd19,  
12'd225,  -12'd166,  12'd154,  12'd167,  12'd118,  -12'd83,  -12'd73,  -12'd177,  12'd29,  -12'd343,  -12'd173,  12'd321,  -12'd4,  -12'd33,  -12'd25,  -12'd291,  
12'd345,  -12'd408,  -12'd209,  12'd28,  -12'd73,  12'd50,  12'd380,  -12'd85,  -12'd37,  12'd376,  12'd26,  12'd37,  12'd12,  12'd721,  12'd58,  -12'd357,  
-12'd458,  12'd255,  12'd256,  -12'd38,  12'd87,  -12'd168,  -12'd230,  12'd8,  12'd23,  12'd258,  12'd67,  -12'd199,  -12'd394,  -12'd64,  12'd82,  -12'd307,  
12'd200,  12'd291,  -12'd74,  -12'd69,  12'd159,  12'd291,  12'd172,  -12'd448,  12'd353,  -12'd116,  12'd167,  12'd265,  -12'd445,  12'd157,  -12'd138,  12'd31,  
-12'd147,  12'd328,  12'd185,  -12'd138,  -12'd223,  12'd384,  -12'd271,  12'd215,  -12'd187,  12'd354,  -12'd305,  12'd66,  12'd242,  12'd161,  -12'd61,  -12'd187,  
12'd335,  -12'd343,  12'd175,  12'd9,  -12'd209,  12'd392,  12'd285,  12'd239,  -12'd444,  12'd27,  -12'd91,  12'd268,  -12'd244,  -12'd44,  -12'd13,  -12'd123,  
12'd263,  12'd201,  12'd493,  12'd133,  12'd324,  12'd9,  12'd286,  12'd31,  -12'd188,  -12'd259,  12'd11,  12'd86,  12'd68,  12'd260,  -12'd111,  -12'd131,  
12'd180,  12'd101,  12'd401,  12'd162,  -12'd96,  -12'd169,  12'd22,  12'd211,  -12'd192,  -12'd413,  12'd167,  12'd164,  12'd28,  12'd134,  12'd36,  -12'd420,  
12'd60,  -12'd75,  12'd34,  -12'd18,  12'd358,  -12'd404,  12'd185,  -12'd87,  -12'd105,  -12'd189,  -12'd198,  -12'd31,  -12'd148,  -12'd4,  12'd262,  12'd147,  
12'd440,  12'd85,  12'd428,  12'd66,  12'd138,  -12'd285,  12'd260,  -12'd74,  -12'd62,  -12'd59,  12'd36,  12'd54,  12'd70,  12'd350,  12'd406,  -12'd18,  
12'd305,  12'd185,  12'd231,  12'd2,  -12'd392,  12'd241,  -12'd59,  12'd119,  -12'd90,  12'd136,  -12'd120,  -12'd101,  -12'd94,  12'd129,  12'd149,  -12'd149,  
-12'd45,  -12'd193,  12'd509,  12'd279,  -12'd92,  -12'd167,  12'd103,  12'd188,  -12'd168,  12'd284,  12'd156,  -12'd391,  -12'd54,  12'd227,  12'd253,  -12'd183,  
12'd348,  12'd141,  12'd513,  12'd106,  -12'd279,  -12'd37,  -12'd84,  12'd89,  -12'd374,  -12'd324,  -12'd397,  -12'd165,  12'd134,  -12'd52,  12'd207,  -12'd64,  
12'd211,  -12'd157,  12'd198,  12'd11,  -12'd247,  12'd136,  -12'd12,  12'd74,  -12'd60,  12'd157,  12'd130,  -12'd7,  -12'd228,  -12'd171,  -12'd123,  -12'd97,  
12'd137,  12'd177,  12'd169,  12'd75,  -12'd123,  -12'd98,  12'd394,  -12'd24,  -12'd123,  -12'd113,  12'd137,  -12'd278,  -12'd381,  12'd380,  12'd283,  12'd347,  
-12'd104,  12'd147,  -12'd94,  -12'd364,  -12'd188,  -12'd24,  12'd57,  -12'd10,  12'd100,  -12'd214,  -12'd192,  -12'd167,  -12'd354,  12'd120,  12'd429,  12'd213,  
12'd263,  -12'd332,  12'd145,  12'd242,  -12'd120,  -12'd96,  -12'd70,  -12'd292,  -12'd321,  12'd218,  -12'd269,  12'd99,  -12'd202,  12'd77,  12'd98,  -12'd15,  
12'd8,  -12'd115,  12'd209,  12'd28,  -12'd171,  12'd262,  12'd35,  12'd85,  12'd188,  -12'd168,  -12'd114,  12'd35,  -12'd139,  12'd73,  -12'd55,  -12'd113,  
-12'd340,  12'd0,  -12'd8,  -12'd134,  -12'd128,  -12'd107,  12'd185,  -12'd241,  -12'd257,  -12'd174,  12'd80,  12'd211,  -12'd151,  -12'd171,  -12'd77,  -12'd453,  
-12'd319,  12'd172,  12'd165,  12'd69,  -12'd176,  12'd191,  12'd190,  -12'd131,  -12'd97,  -12'd216,  -12'd168,  -12'd124,  -12'd34,  12'd307,  12'd258,  12'd114,  
-12'd409,  -12'd236,  12'd226,  12'd12,  -12'd398,  12'd325,  12'd263,  -12'd9,  -12'd194,  12'd53,  12'd271,  12'd156,  12'd22,  12'd2,  12'd124,  -12'd244,  
12'd491,  -12'd573,  12'd519,  12'd255,  -12'd250,  12'd415,  -12'd165,  12'd5,  -12'd10,  -12'd13,  12'd500,  -12'd233,  12'd157,  12'd45,  -12'd125,  12'd174,  
12'd268,  -12'd129,  -12'd396,  12'd116,  -12'd67,  -12'd92,  12'd4,  12'd471,  -12'd166,  12'd66,  -12'd304,  12'd88,  -12'd1,  -12'd283,  -12'd100,  -12'd176,  

-12'd139,  -12'd59,  -12'd42,  -12'd31,  -12'd182,  -12'd117,  -12'd383,  -12'd65,  12'd126,  12'd131,  -12'd48,  12'd36,  12'd53,  12'd289,  12'd108,  -12'd51,  
-12'd253,  -12'd41,  -12'd44,  12'd185,  12'd168,  12'd41,  12'd212,  12'd138,  -12'd28,  -12'd313,  12'd190,  12'd113,  12'd148,  12'd74,  12'd328,  -12'd71,  
-12'd197,  12'd138,  12'd31,  -12'd182,  -12'd270,  12'd15,  12'd141,  -12'd435,  12'd17,  12'd130,  12'd142,  12'd288,  -12'd83,  12'd303,  -12'd57,  -12'd65,  
12'd120,  -12'd260,  -12'd141,  -12'd336,  12'd327,  -12'd69,  12'd22,  12'd199,  12'd192,  -12'd46,  -12'd189,  12'd259,  -12'd55,  -12'd118,  12'd178,  -12'd106,  
-12'd144,  -12'd41,  -12'd137,  -12'd55,  12'd41,  12'd18,  -12'd188,  12'd100,  -12'd275,  12'd200,  -12'd84,  -12'd199,  12'd190,  -12'd248,  12'd0,  12'd167,  
-12'd203,  -12'd106,  -12'd273,  12'd196,  12'd104,  -12'd188,  -12'd100,  -12'd5,  12'd305,  12'd72,  12'd122,  12'd151,  12'd215,  -12'd88,  -12'd123,  -12'd195,  
-12'd295,  -12'd152,  12'd40,  -12'd92,  -12'd9,  -12'd240,  -12'd199,  12'd244,  12'd24,  -12'd208,  12'd19,  -12'd149,  12'd206,  12'd39,  -12'd70,  -12'd93,  
-12'd16,  -12'd173,  -12'd223,  -12'd38,  12'd51,  -12'd148,  -12'd70,  12'd73,  -12'd332,  12'd16,  -12'd227,  -12'd161,  -12'd13,  -12'd303,  -12'd28,  12'd159,  
-12'd179,  -12'd295,  12'd129,  12'd191,  -12'd188,  -12'd66,  -12'd45,  -12'd192,  12'd361,  12'd76,  -12'd68,  -12'd199,  -12'd157,  12'd53,  -12'd6,  12'd0,  
-12'd129,  -12'd150,  -12'd36,  12'd230,  -12'd170,  -12'd104,  12'd324,  -12'd192,  12'd114,  -12'd21,  -12'd61,  -12'd302,  12'd88,  12'd219,  -12'd79,  -12'd44,  
12'd291,  -12'd274,  -12'd368,  12'd106,  -12'd165,  12'd225,  -12'd199,  -12'd250,  12'd264,  -12'd171,  -12'd465,  -12'd224,  -12'd262,  -12'd282,  12'd233,  -12'd114,  
-12'd28,  -12'd427,  12'd111,  12'd181,  12'd268,  -12'd57,  12'd31,  -12'd39,  -12'd230,  12'd283,  12'd182,  -12'd15,  -12'd40,  12'd157,  -12'd24,  -12'd67,  
12'd226,  -12'd141,  -12'd151,  -12'd78,  -12'd113,  12'd18,  -12'd335,  -12'd208,  -12'd191,  -12'd131,  -12'd246,  12'd91,  12'd117,  12'd87,  12'd20,  -12'd48,  
-12'd158,  -12'd303,  12'd77,  -12'd193,  -12'd206,  -12'd378,  -12'd377,  12'd20,  -12'd46,  -12'd166,  12'd302,  -12'd192,  -12'd24,  -12'd183,  -12'd159,  12'd10,  
12'd116,  -12'd80,  -12'd246,  -12'd100,  12'd162,  -12'd272,  12'd198,  12'd11,  -12'd13,  -12'd43,  -12'd78,  -12'd222,  12'd60,  -12'd81,  -12'd75,  12'd21,  
12'd212,  -12'd266,  -12'd253,  -12'd32,  12'd176,  -12'd179,  12'd165,  12'd97,  -12'd11,  12'd285,  -12'd55,  -12'd90,  -12'd142,  -12'd302,  -12'd163,  -12'd70,  
-12'd138,  -12'd74,  -12'd355,  12'd35,  -12'd254,  -12'd150,  -12'd187,  -12'd121,  -12'd89,  -12'd169,  -12'd125,  12'd16,  12'd38,  -12'd219,  -12'd228,  12'd230,  
12'd34,  -12'd116,  12'd120,  -12'd311,  12'd278,  -12'd28,  -12'd424,  -12'd17,  -12'd24,  -12'd399,  -12'd3,  -12'd170,  12'd232,  -12'd187,  -12'd88,  -12'd111,  
12'd23,  12'd177,  12'd246,  -12'd150,  -12'd340,  -12'd263,  -12'd28,  12'd71,  12'd252,  -12'd20,  12'd169,  -12'd130,  12'd150,  12'd302,  -12'd105,  12'd204,  
12'd10,  -12'd331,  12'd164,  12'd134,  -12'd37,  -12'd274,  -12'd136,  12'd362,  -12'd290,  -12'd410,  -12'd242,  12'd64,  -12'd93,  -12'd299,  12'd96,  -12'd47,  
12'd241,  -12'd97,  -12'd257,  -12'd83,  12'd27,  12'd28,  12'd123,  -12'd129,  12'd182,  -12'd9,  12'd22,  12'd33,  12'd95,  -12'd294,  -12'd145,  12'd18,  
12'd119,  12'd137,  -12'd170,  12'd286,  -12'd363,  12'd263,  -12'd66,  -12'd238,  -12'd118,  -12'd96,  -12'd163,  -12'd173,  12'd186,  -12'd40,  12'd143,  12'd158,  
12'd7,  -12'd416,  12'd16,  12'd75,  -12'd120,  -12'd23,  -12'd47,  12'd172,  12'd1,  -12'd156,  12'd267,  -12'd432,  12'd110,  12'd216,  -12'd138,  -12'd131,  
12'd168,  12'd23,  -12'd220,  -12'd100,  12'd208,  -12'd345,  -12'd167,  -12'd137,  12'd196,  -12'd385,  -12'd272,  12'd165,  12'd172,  12'd69,  12'd94,  12'd243,  
-12'd399,  -12'd97,  -12'd374,  12'd11,  -12'd326,  12'd89,  -12'd355,  -12'd96,  12'd218,  -12'd163,  -12'd26,  12'd272,  -12'd45,  -12'd187,  -12'd372,  -12'd92,  

12'd60,  12'd117,  -12'd124,  12'd39,  12'd200,  12'd327,  -12'd121,  -12'd171,  -12'd317,  12'd99,  12'd431,  -12'd210,  12'd371,  -12'd48,  -12'd358,  12'd3,  
-12'd97,  -12'd96,  -12'd416,  12'd454,  -12'd22,  -12'd378,  -12'd651,  12'd0,  12'd202,  12'd37,  -12'd153,  -12'd110,  12'd173,  -12'd797,  12'd104,  12'd100,  
-12'd94,  12'd413,  12'd314,  12'd462,  12'd125,  -12'd23,  -12'd250,  -12'd164,  12'd104,  12'd261,  12'd6,  12'd184,  -12'd279,  -12'd411,  12'd407,  12'd52,  
12'd36,  12'd23,  12'd171,  -12'd130,  -12'd51,  12'd42,  12'd127,  -12'd249,  -12'd66,  12'd62,  -12'd79,  12'd346,  12'd225,  12'd585,  12'd93,  -12'd52,  
-12'd435,  -12'd315,  12'd10,  -12'd44,  12'd36,  -12'd194,  12'd66,  12'd68,  12'd493,  -12'd82,  12'd34,  12'd366,  -12'd410,  -12'd208,  -12'd309,  -12'd250,  
12'd62,  12'd175,  -12'd269,  12'd75,  12'd189,  -12'd193,  -12'd196,  -12'd199,  12'd79,  12'd20,  -12'd24,  -12'd107,  12'd76,  -12'd597,  12'd162,  12'd183,  
-12'd321,  12'd184,  -12'd418,  -12'd200,  12'd381,  12'd115,  12'd252,  -12'd184,  -12'd25,  12'd280,  -12'd58,  12'd112,  -12'd121,  -12'd504,  -12'd57,  -12'd195,  
12'd55,  12'd221,  -12'd18,  -12'd25,  12'd201,  12'd24,  -12'd235,  12'd118,  -12'd513,  -12'd4,  12'd12,  12'd169,  -12'd31,  12'd156,  -12'd343,  12'd572,  
12'd145,  -12'd13,  12'd70,  -12'd421,  12'd157,  12'd385,  12'd477,  -12'd464,  -12'd372,  -12'd146,  -12'd56,  12'd269,  12'd109,  12'd412,  -12'd282,  12'd371,  
12'd9,  12'd24,  12'd12,  -12'd213,  12'd155,  12'd124,  12'd335,  -12'd79,  -12'd282,  -12'd577,  12'd84,  -12'd247,  12'd63,  12'd341,  12'd115,  -12'd272,  
-12'd161,  12'd218,  -12'd374,  -12'd47,  12'd264,  12'd151,  -12'd157,  -12'd29,  12'd456,  -12'd137,  12'd192,  12'd133,  -12'd255,  -12'd201,  12'd31,  12'd202,  
-12'd99,  -12'd122,  -12'd247,  12'd130,  12'd439,  12'd105,  -12'd150,  -12'd237,  12'd62,  12'd260,  -12'd349,  -12'd170,  -12'd44,  -12'd99,  12'd149,  12'd81,  
12'd144,  -12'd90,  12'd154,  -12'd42,  -12'd247,  -12'd73,  -12'd310,  12'd142,  12'd84,  -12'd177,  -12'd127,  12'd173,  12'd309,  -12'd84,  12'd396,  -12'd231,  
12'd161,  12'd79,  12'd189,  12'd235,  -12'd100,  -12'd43,  12'd59,  -12'd347,  12'd275,  12'd26,  12'd164,  12'd298,  12'd239,  12'd11,  -12'd135,  12'd74,  
12'd236,  -12'd81,  12'd57,  12'd287,  12'd219,  -12'd128,  12'd186,  12'd58,  12'd38,  12'd135,  -12'd150,  12'd137,  12'd583,  12'd87,  -12'd315,  12'd57,  
-12'd171,  12'd74,  -12'd424,  -12'd173,  12'd8,  -12'd94,  -12'd59,  -12'd209,  -12'd30,  12'd159,  12'd244,  12'd105,  -12'd62,  -12'd220,  12'd159,  12'd12,  
12'd75,  12'd70,  -12'd11,  -12'd71,  12'd50,  12'd61,  -12'd216,  -12'd367,  12'd588,  -12'd178,  12'd33,  12'd241,  12'd376,  -12'd319,  -12'd109,  -12'd65,  
-12'd216,  12'd374,  12'd252,  -12'd110,  12'd54,  12'd117,  -12'd135,  12'd140,  12'd42,  12'd283,  -12'd9,  -12'd290,  12'd281,  -12'd487,  -12'd151,  12'd384,  
-12'd172,  -12'd277,  -12'd416,  12'd26,  12'd16,  12'd54,  12'd43,  12'd263,  12'd18,  -12'd46,  12'd409,  12'd109,  12'd258,  -12'd330,  -12'd108,  -12'd274,  
-12'd136,  12'd315,  -12'd407,  12'd117,  12'd214,  -12'd387,  -12'd164,  -12'd75,  12'd153,  12'd525,  12'd121,  -12'd76,  12'd223,  -12'd74,  12'd246,  -12'd194,  
-12'd12,  -12'd320,  -12'd122,  -12'd187,  -12'd58,  12'd248,  -12'd229,  -12'd156,  12'd249,  -12'd31,  12'd142,  12'd177,  -12'd62,  -12'd111,  12'd438,  -12'd9,  
12'd218,  12'd209,  12'd161,  -12'd10,  12'd46,  -12'd139,  -12'd245,  12'd96,  12'd53,  -12'd212,  12'd90,  12'd144,  12'd95,  12'd82,  -12'd34,  12'd146,  
12'd67,  -12'd116,  -12'd89,  -12'd10,  12'd318,  12'd82,  -12'd202,  -12'd154,  -12'd153,  12'd274,  -12'd150,  12'd341,  -12'd379,  12'd35,  12'd78,  12'd254,  
-12'd65,  12'd262,  12'd156,  12'd42,  12'd269,  12'd371,  12'd147,  12'd151,  -12'd17,  -12'd138,  -12'd167,  12'd131,  -12'd20,  12'd179,  12'd97,  -12'd119,  
-12'd149,  -12'd196,  12'd88,  12'd207,  12'd26,  -12'd165,  12'd233,  -12'd196,  -12'd6,  12'd449,  -12'd190,  12'd79,  12'd193,  12'd15,  -12'd253,  12'd107,  

12'd210,  -12'd163,  12'd242,  -12'd314,  -12'd403,  -12'd188,  -12'd41,  12'd83,  12'd360,  12'd210,  -12'd83,  12'd300,  -12'd40,  -12'd25,  12'd59,  -12'd218,  
12'd209,  -12'd58,  -12'd190,  12'd176,  -12'd250,  -12'd56,  12'd142,  12'd323,  12'd32,  -12'd277,  -12'd169,  12'd177,  -12'd27,  -12'd58,  -12'd186,  -12'd47,  
-12'd342,  -12'd4,  -12'd184,  12'd93,  12'd62,  12'd109,  12'd87,  -12'd27,  -12'd257,  12'd72,  -12'd259,  12'd326,  -12'd3,  12'd108,  -12'd157,  -12'd179,  
-12'd9,  12'd88,  12'd178,  -12'd389,  -12'd19,  -12'd10,  12'd255,  12'd130,  12'd70,  12'd355,  -12'd125,  12'd358,  -12'd193,  -12'd155,  12'd99,  -12'd152,  
12'd323,  12'd26,  12'd471,  12'd93,  -12'd314,  12'd192,  -12'd321,  12'd274,  -12'd151,  12'd270,  12'd157,  12'd160,  -12'd128,  -12'd170,  12'd245,  12'd375,  
12'd96,  -12'd144,  -12'd14,  -12'd3,  12'd180,  -12'd12,  -12'd252,  12'd432,  12'd466,  12'd380,  -12'd257,  12'd175,  12'd147,  12'd69,  12'd329,  -12'd253,  
-12'd203,  -12'd225,  -12'd19,  12'd204,  -12'd36,  12'd54,  12'd236,  12'd232,  12'd325,  -12'd22,  12'd90,  12'd15,  12'd119,  12'd20,  12'd22,  -12'd24,  
-12'd49,  -12'd186,  12'd93,  12'd57,  -12'd239,  12'd173,  -12'd160,  12'd29,  12'd64,  12'd136,  -12'd63,  12'd169,  12'd327,  -12'd201,  12'd28,  12'd119,  
-12'd210,  12'd253,  12'd163,  -12'd73,  -12'd84,  -12'd175,  12'd46,  12'd145,  12'd62,  -12'd241,  -12'd136,  12'd21,  12'd168,  -12'd88,  12'd36,  12'd182,  
12'd456,  -12'd7,  12'd246,  -12'd1,  12'd134,  -12'd372,  -12'd252,  12'd191,  -12'd155,  12'd55,  12'd171,  12'd93,  12'd472,  12'd15,  -12'd60,  12'd503,  
12'd116,  12'd312,  12'd80,  12'd90,  12'd581,  12'd206,  -12'd143,  12'd395,  -12'd61,  -12'd401,  -12'd144,  -12'd43,  12'd418,  12'd246,  -12'd155,  12'd122,  
-12'd30,  12'd118,  12'd347,  12'd403,  12'd120,  -12'd69,  12'd397,  12'd48,  12'd166,  -12'd485,  12'd128,  -12'd192,  12'd14,  12'd62,  -12'd226,  12'd135,  
-12'd61,  12'd203,  -12'd74,  -12'd66,  -12'd49,  12'd233,  12'd54,  -12'd12,  12'd137,  -12'd410,  12'd194,  12'd113,  -12'd2,  -12'd541,  12'd99,  -12'd90,  
12'd189,  -12'd41,  -12'd289,  12'd84,  -12'd202,  -12'd407,  -12'd261,  12'd54,  -12'd427,  -12'd369,  12'd0,  12'd174,  12'd235,  12'd470,  12'd164,  -12'd269,  
12'd477,  -12'd36,  -12'd28,  12'd284,  -12'd48,  12'd175,  12'd199,  -12'd175,  -12'd253,  -12'd268,  12'd1,  -12'd163,  12'd507,  -12'd219,  -12'd169,  12'd264,  
12'd52,  12'd183,  -12'd236,  -12'd188,  -12'd60,  12'd270,  -12'd143,  -12'd90,  -12'd319,  -12'd245,  -12'd315,  12'd489,  -12'd18,  -12'd42,  -12'd174,  -12'd191,  
-12'd52,  -12'd75,  -12'd130,  -12'd99,  12'd190,  -12'd239,  -12'd207,  -12'd34,  12'd35,  12'd180,  -12'd417,  -12'd11,  -12'd50,  12'd244,  12'd107,  12'd256,  
-12'd377,  12'd325,  -12'd179,  -12'd54,  12'd51,  -12'd26,  12'd42,  -12'd383,  -12'd140,  -12'd164,  12'd171,  12'd10,  -12'd145,  -12'd147,  -12'd29,  12'd122,  
-12'd24,  -12'd139,  -12'd196,  -12'd84,  12'd23,  12'd288,  -12'd230,  12'd35,  -12'd128,  12'd111,  12'd171,  12'd43,  12'd236,  12'd17,  12'd31,  12'd195,  
-12'd196,  -12'd59,  12'd611,  -12'd292,  12'd109,  -12'd96,  12'd8,  12'd128,  -12'd123,  12'd22,  12'd160,  12'd82,  12'd221,  12'd142,  -12'd228,  -12'd193,  
12'd193,  12'd425,  12'd294,  -12'd73,  12'd31,  -12'd62,  -12'd625,  -12'd2,  -12'd415,  12'd214,  -12'd115,  12'd254,  12'd215,  12'd200,  12'd137,  -12'd369,  
12'd5,  -12'd219,  -12'd240,  -12'd48,  -12'd48,  -12'd343,  -12'd481,  -12'd21,  -12'd260,  12'd75,  -12'd282,  -12'd2,  -12'd138,  12'd286,  12'd175,  12'd107,  
-12'd142,  12'd29,  -12'd11,  -12'd108,  12'd67,  -12'd41,  12'd92,  12'd60,  -12'd367,  -12'd503,  -12'd131,  -12'd35,  -12'd145,  -12'd147,  -12'd120,  -12'd193,  
12'd456,  -12'd185,  -12'd141,  -12'd12,  12'd2,  12'd85,  -12'd287,  -12'd182,  -12'd23,  -12'd131,  -12'd69,  12'd337,  12'd25,  12'd428,  12'd114,  -12'd28,  
12'd124,  -12'd37,  12'd256,  12'd292,  12'd149,  -12'd6,  12'd232,  -12'd206,  -12'd111,  -12'd612,  -12'd355,  12'd97,  12'd168,  12'd104,  -12'd194,  -12'd125,  

-12'd252,  12'd16,  12'd110,  12'd95,  12'd172,  12'd175,  -12'd647,  12'd15,  -12'd34,  -12'd52,  -12'd155,  12'd244,  -12'd54,  12'd35,  12'd69,  -12'd79,  
12'd162,  -12'd92,  -12'd11,  -12'd273,  12'd19,  -12'd1,  12'd173,  -12'd55,  12'd142,  -12'd186,  -12'd67,  -12'd57,  12'd340,  -12'd383,  12'd300,  -12'd69,  
-12'd164,  12'd228,  12'd114,  12'd103,  -12'd165,  -12'd177,  -12'd59,  12'd86,  12'd141,  -12'd415,  -12'd346,  -12'd73,  12'd194,  12'd110,  12'd96,  12'd93,  
12'd33,  12'd539,  12'd40,  -12'd241,  12'd207,  12'd56,  -12'd407,  -12'd23,  12'd339,  12'd216,  -12'd428,  -12'd181,  12'd84,  -12'd135,  12'd353,  12'd285,  
12'd339,  -12'd140,  12'd218,  12'd214,  -12'd116,  12'd13,  -12'd409,  12'd175,  12'd123,  12'd256,  -12'd270,  12'd44,  -12'd198,  -12'd225,  -12'd34,  -12'd671,  
-12'd153,  12'd368,  12'd94,  -12'd49,  12'd152,  12'd58,  12'd326,  -12'd205,  12'd12,  -12'd181,  12'd58,  -12'd73,  12'd193,  12'd248,  12'd73,  12'd176,  
12'd96,  -12'd82,  -12'd234,  12'd219,  12'd99,  12'd54,  12'd478,  12'd84,  12'd14,  -12'd227,  12'd324,  12'd48,  12'd17,  -12'd442,  -12'd225,  12'd11,  
-12'd348,  12'd594,  -12'd239,  -12'd14,  12'd207,  12'd21,  12'd161,  12'd111,  -12'd43,  -12'd79,  -12'd168,  12'd107,  12'd41,  12'd69,  -12'd417,  -12'd160,  
-12'd283,  12'd792,  -12'd47,  12'd214,  12'd260,  -12'd308,  -12'd128,  -12'd37,  12'd197,  -12'd73,  12'd4,  12'd329,  12'd66,  -12'd120,  12'd295,  12'd122,  
12'd447,  12'd453,  12'd409,  -12'd190,  12'd279,  12'd160,  12'd32,  -12'd385,  -12'd169,  -12'd76,  12'd64,  12'd153,  12'd136,  -12'd125,  12'd163,  12'd125,  
12'd290,  12'd241,  12'd203,  12'd191,  -12'd114,  12'd187,  12'd70,  12'd70,  -12'd287,  -12'd274,  -12'd238,  12'd362,  12'd214,  12'd99,  -12'd67,  12'd215,  
-12'd97,  -12'd16,  -12'd112,  12'd37,  12'd172,  -12'd133,  12'd200,  12'd106,  12'd462,  -12'd512,  -12'd81,  -12'd135,  -12'd268,  -12'd175,  -12'd90,  12'd60,  
-12'd228,  12'd109,  12'd156,  12'd205,  12'd405,  -12'd424,  12'd39,  12'd158,  -12'd157,  12'd57,  -12'd22,  12'd107,  -12'd324,  12'd93,  -12'd51,  -12'd11,  
12'd256,  -12'd10,  -12'd91,  12'd263,  -12'd385,  12'd258,  -12'd86,  12'd140,  -12'd154,  -12'd221,  12'd92,  12'd162,  -12'd104,  12'd319,  12'd199,  12'd194,  
12'd587,  12'd291,  12'd190,  -12'd18,  -12'd545,  12'd51,  12'd394,  12'd169,  12'd129,  -12'd56,  -12'd80,  12'd203,  -12'd112,  -12'd73,  12'd395,  -12'd283,  
-12'd52,  -12'd96,  -12'd20,  12'd54,  -12'd157,  -12'd99,  12'd315,  12'd7,  -12'd285,  -12'd269,  -12'd56,  -12'd216,  -12'd311,  -12'd111,  12'd24,  -12'd205,  
12'd225,  12'd5,  -12'd391,  12'd345,  12'd58,  12'd97,  12'd196,  -12'd169,  12'd181,  -12'd105,  -12'd369,  -12'd29,  -12'd210,  -12'd281,  12'd357,  12'd36,  
12'd95,  12'd159,  -12'd179,  12'd30,  -12'd68,  12'd213,  12'd322,  -12'd90,  12'd340,  12'd294,  12'd22,  -12'd186,  -12'd79,  -12'd97,  -12'd53,  -12'd412,  
12'd340,  12'd326,  12'd383,  12'd109,  -12'd40,  12'd348,  12'd6,  12'd170,  -12'd77,  12'd179,  12'd85,  -12'd73,  12'd193,  -12'd138,  12'd114,  -12'd29,  
12'd94,  -12'd7,  -12'd93,  12'd110,  12'd44,  12'd98,  -12'd14,  12'd65,  12'd47,  -12'd146,  12'd81,  -12'd215,  12'd331,  -12'd248,  12'd78,  12'd369,  
12'd88,  12'd105,  12'd221,  -12'd100,  -12'd237,  -12'd383,  -12'd394,  -12'd174,  -12'd504,  12'd266,  -12'd681,  12'd59,  -12'd149,  12'd0,  -12'd163,  -12'd355,  
12'd239,  12'd189,  12'd418,  12'd39,  -12'd116,  12'd484,  -12'd11,  -12'd102,  -12'd75,  12'd237,  -12'd155,  -12'd93,  12'd20,  12'd399,  12'd98,  12'd77,  
-12'd191,  -12'd100,  -12'd53,  12'd176,  -12'd55,  12'd42,  -12'd253,  12'd92,  12'd42,  -12'd19,  12'd50,  -12'd141,  12'd240,  -12'd161,  12'd1,  -12'd337,  
-12'd402,  -12'd259,  -12'd234,  -12'd100,  12'd484,  12'd1,  12'd232,  12'd189,  -12'd588,  12'd224,  -12'd339,  -12'd45,  -12'd113,  -12'd174,  12'd331,  12'd145,  
-12'd437,  -12'd102,  -12'd616,  12'd212,  12'd191,  12'd16,  -12'd96,  12'd98,  -12'd331,  -12'd78,  -12'd53,  -12'd258,  -12'd273,  -12'd168,  -12'd176,  12'd18,  

-12'd239,  12'd548,  -12'd211,  -12'd16,  12'd309,  12'd326,  -12'd181,  12'd170,  -12'd433,  -12'd155,  -12'd100,  -12'd40,  12'd227,  -12'd126,  12'd73,  12'd205,  
12'd86,  12'd463,  -12'd232,  -12'd2,  12'd336,  12'd526,  -12'd458,  -12'd273,  -12'd128,  12'd169,  -12'd103,  12'd28,  12'd17,  12'd105,  12'd318,  12'd488,  
-12'd14,  12'd32,  12'd184,  -12'd264,  12'd206,  -12'd148,  12'd522,  12'd12,  -12'd81,  -12'd210,  12'd8,  12'd211,  12'd115,  12'd460,  -12'd240,  -12'd50,  
-12'd254,  -12'd216,  12'd249,  -12'd28,  -12'd433,  -12'd106,  -12'd61,  -12'd195,  12'd314,  12'd22,  12'd237,  12'd11,  -12'd279,  12'd429,  -12'd224,  12'd146,  
-12'd572,  -12'd609,  12'd206,  -12'd30,  -12'd333,  -12'd357,  12'd10,  -12'd258,  -12'd5,  -12'd194,  -12'd98,  -12'd329,  -12'd457,  -12'd194,  12'd101,  -12'd25,  
-12'd8,  -12'd127,  12'd107,  12'd10,  -12'd114,  -12'd113,  -12'd284,  12'd282,  -12'd276,  -12'd16,  12'd172,  12'd159,  12'd244,  -12'd240,  -12'd311,  12'd437,  
12'd313,  12'd655,  -12'd390,  -12'd28,  12'd71,  12'd90,  -12'd140,  12'd211,  12'd147,  -12'd239,  -12'd317,  12'd90,  12'd178,  12'd224,  12'd161,  12'd232,  
12'd110,  12'd34,  -12'd108,  -12'd45,  -12'd228,  -12'd107,  12'd438,  -12'd14,  -12'd115,  -12'd279,  12'd183,  12'd118,  12'd149,  12'd209,  -12'd8,  12'd102,  
12'd235,  12'd41,  12'd451,  -12'd394,  12'd192,  -12'd54,  12'd436,  12'd114,  12'd139,  12'd99,  12'd54,  12'd174,  -12'd479,  12'd421,  -12'd340,  12'd158,  
12'd31,  -12'd13,  12'd398,  12'd29,  -12'd115,  12'd16,  12'd249,  12'd281,  -12'd118,  -12'd144,  -12'd223,  12'd258,  12'd108,  -12'd483,  -12'd334,  -12'd405,  
-12'd231,  12'd162,  -12'd182,  12'd93,  -12'd70,  -12'd252,  -12'd384,  -12'd109,  -12'd144,  -12'd169,  12'd419,  -12'd190,  -12'd230,  12'd25,  12'd25,  12'd42,  
12'd454,  12'd51,  -12'd113,  -12'd77,  -12'd284,  12'd182,  -12'd423,  -12'd2,  -12'd65,  -12'd120,  -12'd359,  12'd370,  -12'd159,  12'd89,  -12'd47,  -12'd246,  
-12'd29,  12'd11,  12'd260,  -12'd247,  -12'd85,  12'd177,  12'd200,  12'd437,  12'd238,  -12'd354,  12'd10,  -12'd195,  -12'd92,  -12'd29,  12'd60,  12'd223,  
-12'd166,  12'd266,  -12'd36,  12'd369,  12'd240,  12'd39,  12'd135,  12'd36,  12'd97,  12'd159,  -12'd165,  -12'd284,  12'd45,  -12'd4,  -12'd201,  -12'd201,  
-12'd19,  -12'd347,  12'd191,  12'd247,  -12'd77,  -12'd13,  -12'd458,  -12'd34,  12'd315,  12'd178,  12'd121,  12'd298,  -12'd109,  -12'd187,  12'd160,  12'd310,  
12'd0,  -12'd15,  12'd258,  12'd263,  -12'd335,  12'd30,  12'd135,  12'd280,  12'd259,  -12'd175,  12'd246,  -12'd305,  -12'd22,  12'd134,  -12'd122,  -12'd229,  
12'd274,  -12'd288,  12'd196,  -12'd69,  12'd241,  12'd39,  12'd492,  -12'd53,  -12'd128,  -12'd380,  12'd320,  -12'd27,  -12'd330,  -12'd191,  12'd112,  12'd204,  
12'd3,  12'd29,  -12'd48,  -12'd253,  -12'd54,  12'd30,  -12'd131,  12'd89,  12'd81,  -12'd183,  -12'd90,  -12'd239,  -12'd74,  -12'd40,  -12'd355,  12'd51,  
12'd26,  -12'd156,  -12'd491,  -12'd1,  -12'd17,  -12'd144,  -12'd569,  12'd79,  12'd216,  12'd172,  -12'd363,  12'd159,  -12'd48,  12'd389,  12'd230,  12'd442,  
12'd246,  12'd146,  12'd301,  12'd158,  12'd196,  12'd417,  12'd200,  -12'd95,  12'd232,  12'd516,  12'd198,  12'd168,  12'd37,  -12'd397,  12'd132,  12'd106,  
12'd180,  -12'd41,  12'd32,  12'd229,  -12'd107,  12'd375,  12'd309,  12'd107,  12'd258,  12'd269,  12'd235,  -12'd39,  12'd132,  -12'd81,  12'd45,  -12'd119,  
12'd183,  -12'd44,  12'd7,  12'd52,  -12'd78,  -12'd275,  -12'd126,  -12'd38,  -12'd18,  -12'd377,  -12'd67,  -12'd382,  12'd195,  12'd86,  -12'd379,  -12'd98,  
-12'd333,  -12'd129,  -12'd171,  -12'd155,  12'd342,  -12'd257,  -12'd232,  -12'd7,  -12'd370,  12'd425,  -12'd82,  12'd230,  12'd281,  -12'd196,  12'd64,  -12'd66,  
12'd62,  12'd151,  -12'd70,  -12'd417,  -12'd158,  12'd49,  -12'd591,  -12'd199,  12'd530,  12'd465,  -12'd207,  12'd160,  -12'd31,  -12'd233,  -12'd230,  12'd11,  
12'd236,  -12'd7,  12'd15,  -12'd106,  -12'd2,  12'd328,  -12'd32,  -12'd5,  12'd114,  12'd91,  12'd26,  12'd240,  12'd488,  -12'd60,  12'd260,  -12'd42,  

-12'd461,  -12'd651,  -12'd327,  -12'd440,  12'd232,  -12'd278,  12'd299,  -12'd255,  -12'd286,  12'd272,  -12'd465,  -12'd52,  -12'd117,  -12'd45,  -12'd543,  -12'd555,  
12'd96,  12'd258,  -12'd36,  -12'd325,  -12'd352,  -12'd256,  -12'd111,  -12'd4,  -12'd511,  -12'd171,  -12'd226,  -12'd148,  -12'd137,  12'd490,  -12'd315,  -12'd259,  
12'd614,  -12'd47,  12'd533,  12'd263,  -12'd243,  12'd178,  12'd269,  -12'd102,  -12'd121,  -12'd411,  -12'd4,  12'd6,  12'd31,  12'd444,  -12'd265,  -12'd261,  
12'd171,  -12'd2,  -12'd75,  12'd142,  -12'd301,  -12'd186,  12'd107,  12'd27,  12'd116,  -12'd47,  12'd350,  12'd223,  -12'd181,  -12'd351,  -12'd14,  -12'd21,  
12'd111,  12'd78,  12'd52,  12'd91,  -12'd132,  -12'd143,  -12'd33,  12'd153,  -12'd305,  12'd200,  -12'd51,  12'd149,  12'd72,  -12'd134,  12'd138,  12'd346,  
-12'd462,  -12'd32,  -12'd674,  -12'd85,  12'd36,  -12'd136,  -12'd219,  12'd11,  12'd238,  12'd62,  12'd11,  -12'd69,  -12'd12,  -12'd339,  -12'd34,  -12'd56,  
12'd167,  12'd147,  12'd195,  12'd198,  12'd202,  -12'd105,  -12'd433,  -12'd367,  -12'd365,  -12'd311,  12'd329,  12'd230,  -12'd40,  12'd521,  -12'd144,  -12'd126,  
12'd344,  -12'd5,  12'd304,  -12'd38,  -12'd365,  -12'd51,  -12'd198,  12'd260,  12'd211,  12'd277,  -12'd223,  12'd87,  -12'd335,  12'd251,  -12'd275,  -12'd77,  
-12'd35,  12'd212,  12'd21,  -12'd178,  12'd116,  12'd113,  12'd144,  12'd57,  -12'd160,  12'd129,  12'd273,  -12'd87,  12'd119,  12'd348,  12'd257,  -12'd12,  
-12'd3,  -12'd416,  -12'd555,  12'd137,  -12'd108,  -12'd471,  12'd119,  -12'd64,  12'd333,  -12'd322,  -12'd18,  -12'd37,  -12'd621,  12'd114,  12'd69,  12'd36,  
-12'd97,  12'd25,  -12'd380,  12'd250,  12'd121,  -12'd260,  -12'd711,  12'd84,  12'd194,  -12'd54,  12'd240,  -12'd79,  -12'd137,  -12'd477,  12'd241,  12'd15,  
-12'd31,  -12'd191,  -12'd12,  -12'd137,  -12'd397,  -12'd617,  -12'd64,  -12'd556,  -12'd196,  12'd190,  -12'd149,  -12'd263,  -12'd35,  12'd449,  -12'd163,  -12'd98,  
12'd264,  -12'd5,  12'd216,  -12'd123,  -12'd108,  -12'd244,  12'd205,  12'd307,  -12'd40,  -12'd53,  -12'd289,  12'd96,  12'd180,  12'd310,  -12'd120,  -12'd9,  
-12'd32,  12'd293,  12'd556,  -12'd200,  -12'd337,  12'd192,  12'd476,  -12'd143,  12'd276,  -12'd375,  -12'd6,  -12'd2,  -12'd278,  12'd91,  -12'd42,  12'd51,  
12'd392,  12'd307,  -12'd299,  12'd111,  -12'd222,  -12'd446,  12'd164,  12'd348,  -12'd31,  -12'd694,  12'd269,  -12'd157,  -12'd203,  -12'd337,  12'd240,  -12'd617,  
-12'd23,  12'd111,  -12'd81,  -12'd64,  12'd347,  12'd71,  -12'd64,  12'd35,  -12'd171,  12'd197,  12'd20,  -12'd752,  -12'd322,  -12'd210,  -12'd127,  -12'd225,  
-12'd19,  -12'd591,  -12'd29,  -12'd235,  12'd191,  -12'd309,  12'd279,  -12'd268,  -12'd860,  12'd261,  12'd81,  12'd41,  12'd277,  12'd30,  12'd303,  -12'd187,  
-12'd6,  -12'd333,  12'd357,  -12'd222,  -12'd647,  -12'd225,  12'd208,  -12'd273,  12'd163,  -12'd194,  -12'd667,  -12'd157,  -12'd130,  12'd382,  -12'd54,  -12'd726,  
12'd52,  12'd52,  12'd586,  12'd303,  -12'd627,  -12'd354,  -12'd150,  12'd22,  -12'd25,  12'd312,  -12'd81,  12'd9,  -12'd382,  -12'd192,  12'd122,  -12'd801,  
12'd79,  12'd161,  -12'd45,  12'd38,  -12'd799,  -12'd487,  -12'd83,  -12'd24,  -12'd448,  12'd299,  -12'd487,  12'd261,  -12'd64,  -12'd64,  -12'd286,  -12'd491,  
12'd54,  12'd2,  -12'd209,  12'd373,  -12'd165,  -12'd25,  12'd101,  12'd298,  12'd71,  -12'd56,  -12'd187,  -12'd239,  -12'd107,  -12'd261,  12'd5,  12'd193,  
12'd408,  12'd8,  12'd172,  12'd263,  -12'd793,  12'd290,  -12'd169,  -12'd20,  12'd381,  12'd475,  -12'd234,  -12'd55,  -12'd142,  -12'd114,  12'd0,  12'd111,  
12'd38,  -12'd205,  12'd96,  12'd122,  12'd198,  -12'd66,  12'd246,  -12'd41,  12'd359,  12'd649,  12'd104,  -12'd12,  -12'd149,  -12'd243,  12'd155,  12'd183,  
-12'd286,  -12'd343,  12'd204,  12'd239,  12'd51,  -12'd417,  -12'd261,  12'd204,  12'd224,  12'd39,  12'd203,  -12'd86,  -12'd33,  12'd113,  12'd157,  12'd451,  
-12'd85,  -12'd281,  -12'd47,  12'd126,  -12'd13,  -12'd460,  12'd54,  12'd44,  -12'd470,  12'd267,  12'd95,  12'd369,  12'd110,  12'd40,  12'd90,  12'd372,  

12'd146,  -12'd83,  -12'd185,  -12'd5,  12'd438,  -12'd289,  12'd261,  -12'd140,  -12'd54,  12'd280,  12'd82,  -12'd25,  -12'd326,  -12'd289,  -12'd140,  12'd212,  
-12'd140,  -12'd36,  -12'd444,  -12'd297,  12'd192,  12'd99,  12'd341,  12'd98,  12'd22,  -12'd109,  -12'd565,  -12'd47,  12'd346,  12'd85,  -12'd36,  -12'd39,  
-12'd9,  -12'd14,  -12'd157,  -12'd348,  -12'd86,  -12'd9,  -12'd75,  12'd0,  -12'd188,  -12'd331,  -12'd315,  12'd277,  12'd36,  12'd183,  12'd153,  12'd158,  
12'd157,  12'd172,  -12'd310,  -12'd173,  -12'd1,  -12'd7,  12'd259,  -12'd154,  12'd321,  -12'd112,  -12'd19,  12'd68,  12'd127,  12'd752,  12'd188,  12'd241,  
-12'd97,  -12'd58,  12'd29,  -12'd101,  12'd67,  12'd120,  12'd54,  12'd176,  -12'd51,  -12'd4,  12'd13,  -12'd184,  -12'd241,  12'd125,  12'd432,  12'd130,  
12'd14,  12'd412,  -12'd153,  -12'd237,  -12'd228,  -12'd125,  12'd346,  -12'd382,  -12'd153,  12'd240,  12'd254,  12'd78,  12'd4,  -12'd516,  -12'd4,  -12'd94,  
12'd236,  12'd241,  -12'd118,  -12'd118,  12'd42,  -12'd77,  -12'd117,  -12'd255,  12'd232,  12'd349,  -12'd73,  -12'd192,  -12'd158,  -12'd218,  -12'd20,  12'd57,  
-12'd43,  12'd310,  12'd23,  -12'd276,  12'd130,  12'd341,  -12'd123,  12'd37,  12'd77,  -12'd73,  12'd119,  -12'd41,  -12'd14,  -12'd21,  -12'd134,  -12'd67,  
12'd222,  12'd0,  12'd334,  12'd181,  12'd137,  12'd119,  12'd247,  12'd25,  -12'd171,  -12'd330,  12'd30,  12'd194,  -12'd81,  12'd78,  -12'd122,  -12'd247,  
12'd10,  12'd225,  12'd315,  12'd304,  -12'd117,  12'd386,  -12'd120,  12'd2,  12'd212,  -12'd144,  12'd75,  -12'd64,  -12'd257,  12'd269,  12'd374,  -12'd365,  
12'd3,  12'd175,  -12'd223,  12'd27,  -12'd342,  12'd117,  12'd198,  -12'd67,  -12'd45,  12'd95,  -12'd297,  12'd489,  12'd120,  -12'd34,  12'd153,  12'd15,  
-12'd39,  -12'd22,  -12'd254,  -12'd114,  -12'd38,  -12'd199,  -12'd72,  12'd23,  12'd540,  12'd56,  -12'd395,  12'd56,  -12'd306,  -12'd3,  -12'd20,  -12'd232,  
12'd103,  12'd191,  -12'd386,  12'd311,  12'd247,  -12'd276,  12'd139,  12'd24,  12'd73,  12'd13,  -12'd50,  12'd105,  -12'd134,  -12'd30,  -12'd145,  12'd200,  
12'd347,  -12'd30,  12'd155,  12'd90,  -12'd277,  12'd163,  12'd21,  12'd220,  12'd144,  12'd225,  -12'd32,  -12'd39,  -12'd111,  12'd126,  12'd360,  12'd77,  
12'd228,  12'd111,  -12'd59,  12'd146,  -12'd49,  12'd308,  12'd144,  12'd218,  -12'd101,  -12'd111,  -12'd109,  12'd23,  12'd334,  12'd49,  12'd109,  12'd161,  
12'd231,  12'd213,  12'd284,  12'd405,  12'd108,  12'd57,  12'd233,  12'd246,  -12'd173,  12'd160,  12'd50,  -12'd178,  12'd165,  12'd264,  12'd304,  -12'd48,  
12'd289,  -12'd105,  12'd308,  12'd80,  -12'd231,  -12'd107,  -12'd63,  12'd57,  -12'd1,  -12'd345,  -12'd87,  -12'd170,  -12'd189,  12'd67,  12'd228,  -12'd287,  
12'd303,  12'd159,  -12'd544,  12'd157,  12'd203,  12'd56,  -12'd280,  12'd283,  -12'd475,  -12'd64,  12'd213,  -12'd85,  12'd344,  -12'd80,  -12'd0,  12'd223,  
12'd78,  -12'd286,  12'd43,  -12'd12,  12'd314,  12'd106,  -12'd290,  12'd317,  -12'd290,  12'd28,  -12'd290,  -12'd162,  12'd85,  12'd316,  -12'd113,  12'd452,  
12'd114,  12'd142,  -12'd13,  12'd415,  12'd88,  12'd241,  12'd232,  12'd77,  12'd106,  12'd206,  12'd126,  12'd47,  12'd280,  12'd229,  -12'd0,  -12'd124,  
12'd183,  -12'd52,  12'd165,  12'd477,  12'd614,  12'd315,  -12'd351,  12'd339,  -12'd372,  12'd104,  12'd24,  12'd41,  12'd380,  12'd62,  12'd405,  12'd32,  
-12'd417,  12'd47,  12'd152,  12'd386,  12'd153,  -12'd29,  -12'd141,  12'd171,  -12'd13,  -12'd62,  -12'd103,  -12'd83,  -12'd130,  12'd377,  12'd198,  -12'd90,  
-12'd237,  12'd313,  -12'd276,  -12'd278,  -12'd156,  -12'd28,  -12'd346,  12'd139,  -12'd566,  -12'd173,  12'd302,  -12'd12,  -12'd79,  -12'd533,  -12'd313,  -12'd96,  
12'd122,  -12'd58,  12'd130,  12'd289,  -12'd121,  12'd256,  12'd76,  12'd357,  12'd89,  12'd105,  -12'd154,  12'd221,  -12'd87,  -12'd232,  -12'd363,  -12'd239,  
12'd64,  12'd2,  12'd110,  12'd127,  -12'd195,  12'd202,  12'd172,  12'd73,  12'd395,  12'd14,  12'd34,  12'd42,  12'd309,  -12'd243,  -12'd82,  -12'd51,  

12'd39,  12'd203,  -12'd172,  -12'd388,  12'd31,  -12'd270,  12'd242,  -12'd484,  -12'd362,  -12'd251,  -12'd195,  12'd293,  -12'd108,  12'd72,  -12'd33,  -12'd349,  
12'd158,  -12'd114,  -12'd64,  -12'd175,  -12'd24,  -12'd4,  12'd24,  -12'd230,  -12'd381,  12'd5,  -12'd78,  12'd33,  -12'd188,  12'd136,  12'd112,  12'd301,  
12'd224,  12'd453,  -12'd222,  -12'd105,  12'd190,  -12'd101,  12'd230,  -12'd280,  -12'd63,  12'd242,  12'd157,  12'd210,  -12'd362,  12'd67,  -12'd11,  12'd100,  
12'd350,  -12'd222,  12'd228,  12'd145,  -12'd219,  -12'd176,  12'd173,  -12'd513,  -12'd124,  12'd323,  12'd147,  -12'd75,  -12'd48,  -12'd47,  12'd211,  12'd123,  
-12'd294,  -12'd669,  -12'd251,  -12'd333,  -12'd46,  12'd28,  12'd186,  12'd63,  -12'd282,  -12'd342,  -12'd143,  12'd153,  12'd77,  -12'd332,  -12'd281,  12'd218,  
-12'd12,  -12'd105,  12'd130,  -12'd429,  -12'd373,  -12'd126,  12'd91,  -12'd334,  12'd258,  -12'd188,  12'd402,  12'd13,  -12'd461,  12'd74,  -12'd188,  12'd97,  
-12'd67,  12'd242,  -12'd44,  -12'd57,  12'd135,  12'd234,  12'd24,  -12'd209,  -12'd333,  -12'd54,  -12'd264,  12'd59,  -12'd5,  12'd57,  -12'd330,  -12'd369,  
12'd108,  -12'd18,  -12'd182,  12'd123,  -12'd244,  12'd39,  12'd197,  -12'd416,  -12'd100,  -12'd4,  -12'd190,  12'd211,  -12'd215,  -12'd28,  12'd6,  12'd347,  
12'd225,  12'd326,  12'd131,  -12'd518,  -12'd202,  12'd85,  12'd413,  12'd159,  -12'd140,  12'd446,  12'd14,  12'd83,  12'd109,  12'd399,  -12'd148,  12'd64,  
12'd182,  12'd296,  12'd528,  -12'd291,  -12'd242,  -12'd324,  12'd88,  -12'd216,  12'd297,  -12'd316,  -12'd65,  -12'd288,  -12'd376,  12'd16,  -12'd271,  12'd155,  
-12'd384,  -12'd264,  12'd363,  12'd203,  -12'd22,  -12'd25,  -12'd102,  12'd147,  12'd190,  12'd227,  -12'd352,  -12'd181,  -12'd258,  -12'd109,  12'd150,  -12'd157,  
12'd20,  12'd109,  -12'd103,  -12'd5,  -12'd325,  12'd77,  12'd233,  12'd129,  -12'd73,  -12'd64,  12'd64,  -12'd196,  12'd120,  -12'd8,  -12'd116,  12'd9,  
12'd370,  12'd90,  12'd575,  -12'd40,  -12'd376,  12'd365,  12'd281,  12'd158,  -12'd171,  -12'd46,  12'd90,  12'd179,  12'd122,  12'd474,  12'd113,  12'd305,  
12'd297,  12'd387,  12'd446,  -12'd50,  -12'd343,  -12'd160,  12'd413,  12'd505,  12'd210,  12'd111,  12'd231,  12'd285,  -12'd85,  12'd386,  12'd108,  -12'd310,  
12'd114,  12'd117,  -12'd199,  -12'd155,  12'd41,  -12'd274,  12'd137,  -12'd19,  -12'd242,  -12'd370,  -12'd221,  -12'd144,  12'd127,  12'd129,  -12'd339,  -12'd171,  
12'd242,  -12'd350,  -12'd158,  -12'd269,  -12'd389,  12'd188,  12'd289,  -12'd100,  12'd377,  -12'd22,  12'd310,  -12'd30,  -12'd79,  12'd133,  -12'd90,  -12'd163,  
12'd59,  12'd167,  12'd70,  12'd142,  -12'd96,  -12'd105,  12'd343,  12'd223,  -12'd229,  -12'd204,  12'd526,  -12'd0,  12'd239,  12'd447,  12'd82,  12'd7,  
-12'd353,  12'd205,  12'd462,  -12'd87,  -12'd199,  12'd99,  12'd402,  12'd114,  12'd158,  12'd176,  -12'd303,  -12'd300,  12'd182,  12'd625,  -12'd148,  -12'd31,  
-12'd64,  -12'd259,  12'd97,  12'd40,  12'd22,  -12'd463,  -12'd116,  -12'd5,  -12'd444,  -12'd405,  -12'd408,  -12'd16,  -12'd157,  12'd140,  -12'd255,  -12'd173,  
12'd39,  12'd7,  12'd298,  12'd278,  -12'd600,  -12'd430,  -12'd383,  -12'd212,  -12'd58,  -12'd93,  -12'd245,  -12'd164,  -12'd35,  12'd398,  -12'd82,  -12'd418,  
-12'd311,  12'd227,  -12'd228,  -12'd330,  12'd159,  -12'd33,  12'd566,  12'd257,  -12'd149,  12'd201,  12'd72,  12'd305,  -12'd137,  -12'd547,  -12'd127,  12'd104,  
-12'd164,  12'd70,  -12'd122,  12'd113,  12'd311,  -12'd283,  12'd257,  -12'd40,  12'd325,  12'd206,  12'd173,  -12'd389,  -12'd198,  12'd289,  -12'd196,  -12'd327,  
-12'd67,  -12'd76,  12'd316,  12'd5,  12'd225,  -12'd30,  12'd333,  12'd271,  12'd393,  12'd384,  -12'd22,  -12'd610,  -12'd157,  12'd334,  12'd171,  -12'd262,  
-12'd512,  -12'd106,  -12'd190,  12'd63,  12'd310,  -12'd184,  -12'd241,  -12'd314,  12'd135,  12'd296,  12'd106,  -12'd146,  12'd63,  12'd200,  12'd47,  -12'd231,  
12'd40,  -12'd187,  12'd845,  12'd83,  12'd280,  12'd43,  -12'd199,  -12'd448,  -12'd237,  12'd1242,  12'd89,  12'd626,  12'd556,  -12'd576,  12'd502,  -12'd185,  

-12'd4,  -12'd60,  12'd344,  12'd154,  12'd104,  12'd161,  -12'd312,  12'd290,  12'd341,  12'd171,  -12'd137,  12'd431,  -12'd199,  12'd109,  -12'd31,  -12'd15,  
-12'd122,  -12'd176,  12'd315,  12'd7,  -12'd81,  -12'd120,  -12'd281,  12'd305,  12'd126,  12'd127,  -12'd273,  -12'd195,  12'd117,  12'd289,  12'd243,  -12'd55,  
12'd266,  -12'd518,  12'd187,  -12'd100,  -12'd60,  -12'd71,  12'd170,  -12'd17,  12'd224,  -12'd13,  -12'd39,  -12'd197,  -12'd199,  12'd537,  -12'd138,  -12'd101,  
-12'd329,  -12'd446,  -12'd292,  -12'd291,  -12'd172,  12'd251,  12'd341,  12'd101,  -12'd30,  12'd117,  12'd39,  -12'd116,  -12'd66,  12'd567,  -12'd180,  -12'd218,  
12'd565,  12'd503,  -12'd62,  -12'd93,  12'd312,  12'd110,  12'd157,  -12'd40,  12'd247,  12'd132,  12'd12,  12'd85,  -12'd137,  -12'd18,  -12'd225,  12'd11,  
-12'd223,  -12'd64,  -12'd30,  12'd334,  12'd620,  12'd237,  -12'd366,  12'd198,  -12'd0,  -12'd10,  12'd16,  12'd140,  12'd198,  12'd494,  -12'd118,  12'd421,  
-12'd442,  12'd382,  12'd109,  12'd66,  -12'd259,  -12'd256,  12'd173,  -12'd43,  -12'd188,  -12'd12,  -12'd336,  12'd65,  12'd154,  -12'd55,  12'd384,  12'd89,  
12'd114,  -12'd124,  12'd100,  12'd163,  -12'd59,  -12'd7,  12'd61,  -12'd16,  12'd25,  -12'd249,  12'd350,  -12'd2,  -12'd182,  12'd81,  -12'd12,  12'd15,  
12'd375,  -12'd196,  12'd213,  12'd188,  -12'd54,  -12'd125,  12'd402,  12'd310,  12'd67,  -12'd69,  12'd4,  -12'd51,  12'd288,  12'd104,  -12'd197,  -12'd253,  
12'd693,  -12'd28,  -12'd412,  -12'd0,  -12'd252,  -12'd161,  12'd31,  -12'd30,  -12'd56,  -12'd377,  12'd101,  -12'd182,  12'd155,  -12'd58,  -12'd222,  12'd205,  
-12'd202,  12'd365,  -12'd434,  -12'd182,  -12'd101,  -12'd46,  -12'd201,  12'd232,  -12'd140,  12'd248,  12'd258,  -12'd0,  12'd260,  12'd77,  12'd37,  12'd7,  
-12'd67,  12'd231,  12'd80,  12'd45,  -12'd145,  12'd105,  12'd112,  -12'd166,  -12'd236,  -12'd317,  12'd194,  -12'd24,  12'd344,  12'd15,  12'd128,  12'd370,  
-12'd157,  -12'd268,  12'd151,  12'd98,  -12'd15,  12'd96,  12'd219,  12'd300,  -12'd92,  -12'd145,  12'd51,  12'd107,  12'd483,  -12'd149,  12'd172,  -12'd26,  
12'd171,  12'd4,  12'd205,  12'd300,  12'd86,  -12'd254,  12'd291,  12'd192,  12'd33,  12'd90,  12'd275,  -12'd76,  12'd195,  -12'd462,  -12'd173,  -12'd230,  
-12'd445,  -12'd142,  -12'd332,  -12'd332,  12'd155,  -12'd40,  12'd135,  12'd1,  -12'd449,  12'd71,  12'd247,  -12'd120,  12'd57,  -12'd341,  -12'd140,  12'd51,  
-12'd41,  12'd134,  -12'd276,  -12'd207,  12'd457,  12'd44,  -12'd126,  12'd92,  12'd181,  12'd82,  12'd475,  12'd86,  -12'd379,  -12'd65,  -12'd322,  -12'd64,  
-12'd104,  12'd218,  -12'd50,  -12'd349,  12'd191,  -12'd38,  12'd603,  -12'd53,  -12'd67,  12'd164,  12'd145,  -12'd73,  12'd102,  -12'd202,  -12'd42,  12'd225,  
-12'd4,  12'd113,  12'd70,  12'd38,  -12'd310,  12'd208,  12'd135,  -12'd70,  12'd369,  12'd159,  -12'd243,  -12'd407,  -12'd10,  12'd85,  -12'd123,  12'd43,  
12'd70,  -12'd235,  12'd57,  12'd157,  -12'd427,  12'd197,  -12'd11,  -12'd62,  12'd54,  12'd146,  12'd468,  12'd27,  -12'd136,  12'd336,  -12'd39,  12'd120,  
-12'd109,  -12'd363,  12'd172,  -12'd28,  12'd159,  12'd20,  12'd36,  12'd55,  12'd116,  -12'd295,  12'd50,  12'd163,  -12'd107,  -12'd48,  -12'd189,  12'd123,  
-12'd255,  -12'd341,  -12'd287,  12'd128,  12'd87,  -12'd44,  -12'd64,  -12'd137,  12'd299,  12'd52,  -12'd31,  -12'd106,  12'd101,  -12'd414,  12'd27,  -12'd20,  
-12'd203,  -12'd64,  -12'd125,  -12'd152,  -12'd215,  -12'd137,  12'd277,  12'd267,  12'd539,  12'd179,  12'd192,  12'd62,  12'd38,  12'd382,  -12'd162,  12'd343,  
12'd422,  12'd66,  12'd181,  12'd235,  12'd91,  -12'd191,  12'd403,  -12'd129,  12'd56,  12'd513,  -12'd75,  12'd57,  -12'd149,  12'd599,  12'd69,  12'd39,  
12'd335,  12'd81,  12'd147,  -12'd149,  12'd2,  12'd110,  -12'd35,  -12'd135,  -12'd210,  -12'd37,  12'd221,  -12'd75,  -12'd116,  12'd189,  12'd44,  12'd93,  
12'd380,  -12'd80,  12'd186,  12'd279,  -12'd17,  12'd11,  12'd172,  12'd78,  -12'd503,  -12'd577,  12'd174,  -12'd115,  -12'd35,  12'd201,  -12'd83,  12'd114,  

12'd334,  12'd68,  12'd200,  -12'd22,  12'd60,  -12'd65,  -12'd340,  12'd6,  12'd139,  12'd263,  -12'd494,  12'd90,  -12'd132,  -12'd374,  12'd302,  12'd497,  
-12'd31,  12'd139,  12'd623,  12'd59,  12'd100,  -12'd238,  12'd204,  12'd438,  -12'd542,  12'd114,  -12'd444,  -12'd7,  -12'd689,  12'd403,  -12'd307,  12'd2,  
-12'd183,  -12'd480,  12'd316,  -12'd285,  -12'd437,  -12'd194,  12'd419,  12'd163,  12'd36,  12'd16,  -12'd450,  -12'd76,  -12'd278,  12'd497,  12'd81,  -12'd580,  
-12'd501,  12'd344,  12'd180,  -12'd208,  -12'd503,  -12'd129,  12'd223,  -12'd29,  12'd68,  12'd65,  -12'd8,  -12'd277,  -12'd355,  -12'd180,  -12'd328,  -12'd675,  
-12'd348,  12'd55,  -12'd207,  -12'd241,  -12'd509,  -12'd391,  -12'd443,  -12'd341,  -12'd400,  -12'd134,  -12'd227,  -12'd311,  -12'd630,  -12'd469,  12'd82,  -12'd310,  
-12'd210,  -12'd156,  -12'd403,  12'd258,  12'd215,  12'd393,  12'd270,  -12'd141,  -12'd165,  -12'd140,  -12'd106,  12'd165,  12'd214,  -12'd20,  -12'd377,  -12'd7,  
12'd194,  12'd284,  12'd812,  12'd30,  12'd0,  12'd479,  12'd565,  12'd459,  -12'd215,  12'd78,  -12'd90,  12'd266,  12'd82,  12'd402,  12'd94,  -12'd21,  
-12'd651,  12'd368,  12'd64,  12'd56,  -12'd242,  12'd295,  12'd501,  12'd575,  12'd84,  12'd395,  -12'd89,  -12'd375,  12'd251,  -12'd68,  -12'd64,  -12'd596,  
12'd351,  -12'd382,  12'd327,  -12'd20,  -12'd69,  -12'd314,  -12'd474,  -12'd123,  -12'd91,  12'd440,  -12'd258,  12'd228,  12'd149,  12'd10,  12'd132,  12'd77,  
12'd317,  12'd27,  12'd69,  -12'd135,  12'd181,  12'd203,  -12'd227,  -12'd313,  12'd24,  12'd401,  -12'd527,  12'd344,  -12'd399,  -12'd334,  12'd60,  -12'd126,  
-12'd208,  12'd89,  -12'd26,  12'd50,  12'd252,  12'd274,  12'd254,  -12'd302,  12'd10,  12'd87,  12'd31,  12'd169,  12'd51,  12'd278,  12'd198,  12'd321,  
-12'd351,  12'd18,  -12'd83,  -12'd437,  12'd200,  -12'd27,  12'd735,  -12'd141,  -12'd250,  -12'd117,  -12'd148,  -12'd178,  -12'd91,  12'd192,  12'd318,  -12'd288,  
-12'd170,  12'd255,  12'd115,  12'd395,  12'd97,  -12'd41,  -12'd101,  -12'd285,  12'd202,  -12'd305,  12'd411,  -12'd69,  12'd98,  12'd123,  12'd52,  12'd259,  
12'd115,  12'd183,  12'd310,  -12'd1,  12'd19,  -12'd211,  -12'd220,  -12'd182,  12'd17,  12'd165,  12'd255,  -12'd295,  12'd152,  12'd270,  12'd338,  -12'd31,  
12'd74,  -12'd215,  12'd136,  12'd301,  12'd108,  -12'd187,  12'd221,  -12'd226,  12'd49,  -12'd77,  12'd94,  12'd22,  12'd248,  -12'd423,  12'd169,  12'd86,  
-12'd151,  -12'd25,  12'd241,  -12'd228,  -12'd175,  12'd83,  12'd316,  12'd181,  12'd93,  -12'd118,  12'd275,  -12'd183,  -12'd119,  -12'd148,  12'd51,  -12'd343,  
-12'd223,  -12'd1,  12'd24,  -12'd155,  12'd357,  12'd40,  12'd84,  -12'd222,  -12'd277,  12'd82,  -12'd340,  12'd226,  -12'd156,  -12'd67,  12'd62,  12'd170,  
12'd123,  -12'd18,  12'd273,  -12'd407,  12'd221,  12'd0,  12'd101,  -12'd131,  12'd163,  -12'd15,  -12'd420,  12'd78,  -12'd416,  12'd405,  12'd456,  12'd45,  
12'd575,  -12'd250,  12'd323,  -12'd167,  -12'd343,  -12'd238,  -12'd52,  -12'd311,  12'd249,  12'd211,  12'd53,  12'd217,  -12'd13,  12'd106,  12'd228,  12'd162,  
12'd88,  12'd407,  12'd569,  12'd158,  -12'd1,  12'd500,  12'd166,  -12'd123,  12'd422,  12'd81,  -12'd202,  12'd83,  12'd108,  12'd86,  -12'd64,  -12'd94,  
12'd139,  -12'd270,  12'd183,  -12'd749,  -12'd200,  -12'd424,  -12'd43,  -12'd62,  -12'd505,  -12'd13,  -12'd392,  -12'd191,  -12'd341,  -12'd20,  -12'd149,  -12'd373,  
-12'd41,  12'd55,  -12'd333,  -12'd314,  -12'd105,  -12'd194,  -12'd203,  -12'd244,  -12'd203,  -12'd132,  -12'd530,  -12'd48,  -12'd368,  -12'd239,  -12'd70,  -12'd419,  
12'd423,  -12'd165,  12'd173,  -12'd376,  -12'd478,  12'd418,  12'd17,  12'd149,  -12'd172,  -12'd274,  -12'd212,  -12'd298,  12'd89,  12'd317,  12'd203,  12'd74,  
12'd181,  12'd136,  12'd163,  -12'd27,  -12'd132,  -12'd3,  12'd158,  12'd376,  -12'd290,  -12'd68,  -12'd210,  -12'd161,  -12'd219,  12'd38,  12'd485,  -12'd130,  
-12'd161,  12'd174,  12'd128,  -12'd206,  12'd246,  12'd187,  12'd237,  12'd646,  -12'd118,  12'd19,  -12'd329,  -12'd324,  12'd3,  12'd305,  -12'd24,  12'd202,  

12'd5,  12'd77,  12'd120,  -12'd129,  -12'd338,  -12'd151,  -12'd242,  12'd50,  -12'd382,  12'd221,  -12'd43,  12'd314,  12'd215,  12'd156,  -12'd27,  -12'd77,  
-12'd147,  -12'd29,  -12'd313,  -12'd151,  12'd161,  12'd291,  -12'd101,  -12'd62,  -12'd166,  -12'd293,  12'd352,  12'd184,  -12'd251,  -12'd329,  -12'd392,  12'd163,  
-12'd10,  -12'd118,  -12'd149,  12'd304,  -12'd269,  -12'd130,  12'd88,  12'd288,  12'd11,  12'd101,  -12'd15,  -12'd29,  -12'd1,  12'd95,  12'd330,  -12'd53,  
-12'd26,  -12'd147,  12'd118,  -12'd352,  12'd39,  12'd213,  -12'd151,  12'd81,  -12'd83,  -12'd183,  12'd240,  12'd12,  12'd106,  -12'd359,  12'd147,  -12'd320,  
-12'd89,  -12'd136,  -12'd352,  -12'd325,  -12'd1,  -12'd141,  12'd151,  12'd81,  -12'd156,  -12'd456,  12'd119,  12'd51,  -12'd235,  -12'd315,  12'd185,  -12'd131,  
-12'd76,  -12'd202,  12'd71,  12'd236,  -12'd126,  -12'd47,  -12'd156,  -12'd287,  -12'd61,  -12'd178,  -12'd339,  -12'd86,  12'd135,  -12'd168,  12'd22,  12'd25,  
12'd92,  12'd336,  12'd151,  -12'd237,  -12'd243,  12'd299,  12'd22,  -12'd97,  -12'd271,  12'd248,  -12'd137,  -12'd75,  -12'd299,  12'd266,  12'd21,  12'd97,  
12'd235,  12'd226,  -12'd349,  12'd10,  12'd73,  -12'd92,  -12'd143,  -12'd139,  -12'd117,  12'd65,  -12'd298,  -12'd277,  -12'd8,  -12'd277,  -12'd238,  12'd238,  
12'd28,  12'd131,  12'd118,  -12'd320,  -12'd132,  -12'd105,  12'd223,  -12'd113,  12'd246,  -12'd450,  -12'd55,  -12'd79,  12'd10,  -12'd121,  -12'd31,  -12'd409,  
-12'd49,  -12'd1,  12'd376,  12'd66,  -12'd94,  -12'd275,  -12'd196,  -12'd139,  -12'd32,  12'd16,  -12'd116,  12'd169,  12'd24,  12'd157,  12'd206,  12'd134,  
12'd126,  12'd141,  12'd265,  12'd65,  12'd31,  -12'd118,  12'd146,  12'd194,  -12'd300,  -12'd210,  12'd108,  12'd271,  -12'd340,  -12'd375,  12'd144,  -12'd307,  
12'd160,  12'd63,  -12'd158,  -12'd266,  -12'd148,  12'd224,  -12'd156,  -12'd200,  -12'd22,  12'd111,  -12'd30,  12'd101,  12'd184,  -12'd409,  -12'd69,  -12'd103,  
-12'd179,  12'd114,  -12'd126,  -12'd98,  12'd54,  -12'd165,  12'd57,  -12'd193,  12'd31,  -12'd169,  -12'd223,  -12'd347,  -12'd370,  12'd171,  -12'd19,  12'd56,  
-12'd85,  -12'd376,  -12'd42,  -12'd132,  -12'd209,  -12'd241,  -12'd60,  -12'd41,  -12'd20,  -12'd107,  12'd28,  12'd23,  12'd90,  -12'd154,  -12'd118,  12'd169,  
-12'd26,  -12'd156,  -12'd259,  -12'd3,  -12'd55,  -12'd324,  -12'd157,  12'd65,  -12'd54,  12'd70,  -12'd3,  -12'd340,  12'd85,  -12'd144,  -12'd58,  12'd199,  
-12'd218,  12'd88,  -12'd188,  12'd330,  -12'd9,  -12'd205,  -12'd71,  -12'd81,  -12'd133,  12'd40,  12'd114,  -12'd31,  -12'd366,  -12'd202,  -12'd89,  12'd286,  
12'd18,  -12'd104,  -12'd178,  -12'd294,  -12'd119,  -12'd183,  12'd43,  -12'd118,  -12'd53,  -12'd89,  -12'd19,  -12'd245,  12'd65,  12'd113,  -12'd185,  -12'd203,  
-12'd298,  12'd81,  12'd79,  12'd222,  -12'd1,  -12'd93,  -12'd343,  12'd46,  12'd118,  12'd199,  -12'd380,  -12'd421,  -12'd272,  12'd168,  -12'd181,  -12'd135,  
-12'd266,  -12'd87,  12'd235,  -12'd112,  12'd80,  12'd10,  12'd189,  -12'd155,  -12'd196,  -12'd132,  -12'd58,  -12'd337,  -12'd214,  -12'd210,  12'd2,  12'd111,  
12'd35,  12'd46,  -12'd181,  -12'd238,  -12'd68,  12'd310,  -12'd62,  -12'd105,  12'd162,  -12'd322,  12'd26,  -12'd162,  12'd31,  -12'd103,  12'd186,  -12'd82,  
-12'd387,  12'd21,  12'd82,  -12'd238,  -12'd120,  12'd204,  -12'd6,  12'd111,  -12'd192,  -12'd205,  -12'd302,  12'd29,  -12'd198,  -12'd32,  -12'd196,  12'd1,  
-12'd410,  12'd366,  -12'd104,  -12'd216,  -12'd115,  12'd207,  12'd62,  -12'd167,  -12'd27,  -12'd62,  12'd67,  -12'd3,  -12'd241,  -12'd44,  -12'd125,  -12'd117,  
12'd158,  -12'd166,  12'd43,  -12'd74,  12'd24,  -12'd24,  -12'd48,  -12'd79,  -12'd136,  12'd28,  12'd55,  -12'd220,  -12'd406,  -12'd22,  -12'd81,  -12'd266,  
-12'd176,  -12'd72,  12'd11,  -12'd193,  -12'd39,  12'd96,  12'd74,  -12'd80,  12'd316,  -12'd35,  -12'd189,  12'd345,  12'd66,  12'd32,  -12'd223,  -12'd213,  
-12'd50,  12'd243,  12'd180,  -12'd110,  -12'd29,  12'd28,  -12'd149,  12'd150,  -12'd103,  -12'd207,  -12'd306,  12'd199,  -12'd380,  -12'd438,  -12'd104,  -12'd23,  

-12'd23,  12'd106,  -12'd314,  12'd158,  -12'd415,  -12'd181,  -12'd283,  -12'd220,  12'd37,  -12'd218,  12'd321,  12'd39,  -12'd195,  -12'd415,  -12'd203,  -12'd302,  
-12'd62,  -12'd354,  -12'd219,  12'd50,  -12'd5,  -12'd298,  -12'd324,  12'd294,  12'd239,  12'd167,  -12'd24,  12'd123,  -12'd302,  -12'd374,  12'd136,  -12'd85,  
12'd93,  -12'd342,  -12'd102,  12'd47,  -12'd90,  12'd7,  -12'd487,  -12'd137,  -12'd296,  12'd526,  12'd187,  -12'd219,  12'd183,  -12'd930,  -12'd68,  12'd10,  
-12'd301,  -12'd808,  -12'd307,  12'd392,  12'd248,  12'd229,  -12'd309,  12'd92,  12'd367,  12'd318,  -12'd199,  -12'd164,  -12'd51,  -12'd491,  -12'd263,  12'd67,  
-12'd766,  -12'd419,  12'd167,  12'd84,  -12'd19,  12'd83,  12'd36,  12'd126,  -12'd193,  12'd7,  -12'd384,  -12'd326,  12'd156,  -12'd108,  12'd50,  -12'd605,  
12'd95,  12'd70,  12'd7,  12'd71,  -12'd55,  12'd396,  12'd60,  12'd36,  -12'd77,  -12'd134,  12'd268,  12'd2,  -12'd468,  -12'd148,  -12'd175,  12'd172,  
12'd299,  12'd425,  -12'd37,  12'd78,  -12'd11,  -12'd232,  12'd23,  -12'd46,  12'd265,  12'd28,  -12'd215,  -12'd7,  12'd83,  -12'd341,  -12'd106,  12'd242,  
12'd39,  -12'd97,  -12'd439,  -12'd241,  -12'd85,  12'd419,  -12'd25,  -12'd304,  -12'd41,  -12'd100,  12'd39,  12'd289,  12'd91,  -12'd174,  12'd87,  -12'd0,  
-12'd151,  12'd317,  12'd171,  12'd383,  -12'd181,  -12'd207,  12'd184,  12'd263,  12'd545,  12'd464,  12'd178,  12'd144,  12'd15,  12'd37,  12'd27,  -12'd9,  
-12'd679,  -12'd471,  -12'd298,  12'd62,  -12'd197,  -12'd278,  12'd135,  12'd16,  12'd191,  -12'd373,  12'd137,  -12'd283,  -12'd241,  12'd35,  -12'd157,  -12'd153,  
12'd0,  12'd77,  -12'd4,  -12'd48,  12'd12,  12'd359,  12'd232,  12'd198,  -12'd37,  12'd123,  -12'd465,  12'd38,  12'd268,  12'd217,  -12'd4,  -12'd33,  
-12'd115,  12'd44,  12'd171,  12'd39,  -12'd174,  -12'd174,  12'd65,  12'd119,  12'd64,  -12'd141,  -12'd87,  12'd217,  12'd88,  -12'd316,  12'd161,  -12'd106,  
-12'd86,  12'd245,  -12'd106,  -12'd164,  12'd50,  -12'd287,  -12'd265,  -12'd169,  -12'd346,  12'd60,  12'd215,  -12'd133,  12'd172,  -12'd301,  -12'd35,  12'd150,  
12'd455,  -12'd89,  -12'd20,  -12'd99,  12'd224,  12'd273,  12'd121,  -12'd134,  -12'd65,  -12'd330,  12'd300,  12'd143,  -12'd226,  12'd163,  -12'd50,  12'd72,  
12'd205,  -12'd177,  12'd285,  -12'd25,  12'd123,  -12'd10,  12'd239,  12'd345,  12'd129,  -12'd459,  12'd210,  12'd333,  12'd31,  12'd287,  12'd89,  12'd35,  
12'd75,  -12'd26,  12'd72,  -12'd94,  12'd373,  12'd231,  -12'd115,  12'd4,  -12'd219,  -12'd46,  -12'd152,  12'd112,  12'd43,  12'd395,  -12'd6,  -12'd285,  
12'd19,  -12'd43,  -12'd345,  -12'd17,  -12'd92,  -12'd99,  -12'd265,  12'd276,  12'd2,  -12'd431,  12'd207,  -12'd274,  12'd3,  12'd130,  12'd128,  12'd287,  
-12'd263,  12'd333,  -12'd75,  -12'd257,  12'd48,  -12'd33,  12'd40,  12'd290,  -12'd193,  12'd14,  12'd268,  -12'd128,  -12'd231,  12'd98,  -12'd351,  12'd104,  
12'd397,  12'd394,  12'd205,  -12'd255,  -12'd281,  12'd86,  -12'd15,  -12'd240,  -12'd152,  12'd209,  12'd133,  12'd79,  12'd156,  12'd104,  12'd209,  -12'd173,  
12'd174,  12'd335,  -12'd340,  12'd18,  12'd112,  12'd95,  -12'd116,  12'd246,  -12'd331,  -12'd219,  -12'd134,  -12'd299,  -12'd8,  -12'd39,  12'd259,  12'd68,  
-12'd24,  12'd287,  -12'd47,  -12'd205,  12'd143,  -12'd128,  -12'd323,  -12'd365,  12'd155,  12'd156,  -12'd12,  12'd3,  -12'd457,  -12'd95,  -12'd31,  -12'd165,  
-12'd255,  -12'd397,  12'd327,  12'd81,  -12'd74,  -12'd203,  12'd114,  -12'd125,  12'd168,  12'd61,  12'd70,  -12'd36,  -12'd369,  -12'd210,  -12'd20,  -12'd3,  
-12'd345,  -12'd96,  12'd146,  -12'd140,  12'd43,  12'd196,  12'd373,  -12'd268,  12'd515,  12'd409,  -12'd126,  -12'd195,  -12'd296,  12'd538,  12'd173,  12'd61,  
-12'd190,  -12'd79,  -12'd145,  -12'd349,  12'd39,  12'd273,  -12'd300,  12'd41,  12'd140,  12'd119,  12'd37,  12'd1,  12'd133,  12'd198,  12'd58,  -12'd282,  
-12'd263,  -12'd249,  12'd92,  12'd319,  -12'd405,  -12'd47,  -12'd204,  12'd10,  12'd33,  12'd84,  -12'd253,  -12'd126,  12'd26,  -12'd448,  12'd200,  -12'd278,  

-12'd60,  -12'd17,  -12'd269,  12'd105,  12'd81,  -12'd141,  -12'd55,  12'd104,  -12'd305,  -12'd238,  -12'd308,  12'd117,  -12'd116,  12'd33,  12'd118,  -12'd514,  
12'd42,  12'd360,  -12'd279,  -12'd128,  12'd354,  -12'd6,  -12'd322,  -12'd138,  12'd104,  12'd133,  -12'd159,  12'd133,  -12'd100,  -12'd245,  12'd61,  -12'd90,  
-12'd94,  12'd313,  -12'd376,  -12'd99,  12'd159,  12'd109,  12'd380,  -12'd141,  -12'd291,  12'd148,  12'd131,  12'd218,  -12'd45,  -12'd280,  -12'd126,  12'd148,  
-12'd349,  -12'd94,  12'd143,  -12'd300,  12'd322,  -12'd309,  12'd34,  -12'd344,  12'd183,  -12'd207,  -12'd347,  12'd329,  12'd71,  12'd180,  -12'd191,  12'd274,  
-12'd299,  -12'd481,  -12'd172,  -12'd299,  -12'd205,  -12'd45,  -12'd182,  -12'd64,  -12'd24,  -12'd223,  -12'd87,  -12'd354,  -12'd142,  12'd66,  -12'd252,  -12'd116,  
12'd63,  12'd80,  -12'd42,  12'd208,  -12'd53,  12'd54,  12'd17,  -12'd51,  12'd412,  -12'd121,  -12'd29,  12'd54,  12'd113,  12'd213,  -12'd261,  -12'd195,  
12'd220,  12'd1,  -12'd76,  -12'd253,  -12'd312,  12'd67,  -12'd110,  12'd197,  -12'd253,  -12'd114,  -12'd182,  -12'd135,  12'd239,  -12'd119,  -12'd213,  12'd263,  
12'd389,  -12'd0,  -12'd47,  -12'd66,  -12'd236,  -12'd133,  12'd127,  12'd387,  -12'd188,  -12'd132,  -12'd209,  12'd281,  12'd226,  12'd129,  12'd409,  12'd61,  
-12'd8,  -12'd46,  12'd28,  -12'd65,  12'd10,  12'd87,  12'd533,  -12'd204,  12'd102,  -12'd130,  -12'd12,  12'd481,  12'd97,  12'd704,  12'd59,  -12'd107,  
-12'd288,  12'd10,  -12'd135,  -12'd111,  12'd58,  12'd65,  12'd219,  12'd236,  -12'd99,  12'd148,  -12'd32,  -12'd404,  -12'd57,  12'd165,  -12'd151,  -12'd443,  
-12'd44,  -12'd2,  -12'd84,  -12'd49,  12'd358,  12'd76,  -12'd63,  -12'd122,  -12'd59,  12'd74,  -12'd450,  -12'd114,  -12'd308,  12'd285,  -12'd283,  -12'd133,  
12'd154,  12'd57,  12'd452,  12'd221,  12'd310,  -12'd22,  -12'd274,  -12'd164,  -12'd100,  -12'd350,  12'd58,  12'd285,  12'd39,  -12'd215,  12'd107,  -12'd114,  
12'd117,  12'd138,  12'd99,  -12'd257,  -12'd353,  12'd409,  -12'd208,  12'd353,  12'd119,  -12'd234,  12'd468,  12'd108,  12'd135,  12'd98,  -12'd288,  12'd354,  
-12'd276,  -12'd1,  12'd222,  12'd296,  -12'd349,  -12'd169,  12'd182,  12'd94,  12'd196,  -12'd117,  12'd182,  -12'd146,  12'd119,  12'd195,  12'd181,  -12'd143,  
12'd126,  -12'd223,  -12'd21,  12'd8,  12'd36,  -12'd264,  -12'd198,  -12'd107,  12'd130,  -12'd299,  -12'd19,  -12'd488,  12'd224,  12'd245,  -12'd131,  -12'd356,  
-12'd205,  -12'd102,  -12'd352,  12'd69,  -12'd320,  12'd194,  -12'd84,  -12'd181,  -12'd63,  12'd161,  -12'd83,  -12'd336,  -12'd61,  12'd19,  -12'd262,  12'd137,  
-12'd44,  12'd27,  -12'd195,  12'd225,  -12'd68,  -12'd33,  -12'd185,  12'd363,  12'd154,  -12'd337,  12'd443,  -12'd218,  12'd35,  12'd5,  12'd49,  12'd15,  
12'd137,  -12'd97,  12'd396,  -12'd104,  12'd298,  -12'd287,  -12'd117,  -12'd58,  12'd333,  12'd358,  12'd159,  12'd108,  12'd198,  -12'd16,  -12'd406,  -12'd133,  
12'd233,  -12'd124,  12'd57,  -12'd82,  -12'd256,  12'd121,  -12'd7,  12'd113,  12'd234,  12'd7,  12'd64,  -12'd106,  -12'd93,  12'd318,  12'd32,  -12'd343,  
12'd152,  -12'd350,  -12'd548,  -12'd310,  -12'd298,  -12'd287,  -12'd73,  -12'd295,  -12'd466,  12'd337,  -12'd195,  -12'd88,  12'd43,  12'd113,  -12'd31,  -12'd395,  
12'd53,  12'd15,  12'd29,  -12'd109,  12'd284,  -12'd93,  12'd299,  -12'd351,  -12'd388,  12'd199,  12'd342,  12'd119,  -12'd214,  12'd167,  -12'd9,  12'd304,  
-12'd42,  12'd51,  -12'd202,  12'd108,  12'd44,  -12'd173,  12'd365,  -12'd7,  12'd541,  -12'd0,  12'd169,  -12'd223,  -12'd377,  -12'd65,  12'd41,  12'd237,  
-12'd64,  12'd50,  12'd191,  -12'd113,  12'd217,  -12'd150,  -12'd346,  -12'd61,  12'd52,  -12'd270,  -12'd464,  -12'd67,  12'd64,  12'd532,  12'd59,  12'd64,  
-12'd97,  12'd37,  -12'd37,  12'd103,  -12'd139,  12'd169,  -12'd267,  -12'd228,  -12'd80,  12'd283,  -12'd29,  -12'd32,  -12'd376,  -12'd10,  12'd394,  12'd329,  
-12'd479,  12'd104,  12'd340,  12'd40,  12'd34,  12'd363,  12'd281,  -12'd356,  12'd23,  12'd732,  12'd249,  -12'd321,  -12'd73,  -12'd292,  12'd189,  -12'd148,  

-12'd371,  12'd205,  -12'd100,  12'd315,  -12'd51,  12'd107,  -12'd45,  -12'd241,  12'd236,  -12'd5,  12'd53,  12'd236,  12'd100,  12'd76,  12'd20,  12'd28,  
-12'd190,  12'd307,  12'd48,  12'd343,  -12'd36,  -12'd48,  -12'd203,  12'd414,  -12'd331,  12'd52,  -12'd205,  12'd341,  -12'd74,  12'd250,  -12'd95,  12'd229,  
-12'd189,  -12'd448,  12'd371,  -12'd260,  12'd82,  12'd53,  12'd153,  -12'd116,  12'd437,  12'd22,  -12'd90,  -12'd282,  12'd190,  12'd593,  12'd133,  -12'd87,  
-12'd192,  -12'd454,  -12'd274,  12'd8,  -12'd228,  12'd88,  12'd79,  -12'd16,  -12'd227,  -12'd34,  12'd248,  12'd326,  -12'd204,  -12'd271,  -12'd117,  -12'd138,  
-12'd132,  -12'd287,  -12'd240,  -12'd70,  -12'd184,  -12'd42,  12'd383,  -12'd34,  -12'd342,  -12'd388,  12'd27,  -12'd134,  -12'd95,  12'd164,  12'd10,  12'd109,  
-12'd198,  12'd128,  -12'd137,  -12'd158,  -12'd165,  12'd20,  -12'd185,  12'd16,  -12'd393,  -12'd153,  12'd178,  12'd23,  12'd146,  12'd342,  -12'd64,  12'd30,  
12'd234,  -12'd271,  12'd131,  12'd16,  -12'd43,  -12'd116,  12'd108,  -12'd175,  -12'd312,  -12'd11,  -12'd9,  12'd45,  -12'd269,  -12'd25,  12'd95,  12'd200,  
12'd11,  -12'd344,  -12'd69,  12'd14,  -12'd132,  -12'd131,  -12'd67,  12'd255,  12'd318,  -12'd246,  12'd70,  -12'd56,  -12'd4,  -12'd55,  12'd261,  12'd211,  
-12'd94,  -12'd457,  12'd1,  12'd62,  -12'd242,  -12'd80,  -12'd34,  12'd134,  -12'd54,  -12'd51,  12'd11,  -12'd86,  -12'd36,  -12'd54,  12'd94,  -12'd317,  
-12'd292,  12'd83,  -12'd370,  -12'd60,  -12'd456,  12'd403,  -12'd215,  12'd98,  12'd130,  -12'd162,  12'd159,  -12'd153,  12'd120,  -12'd31,  -12'd75,  12'd356,  
-12'd141,  -12'd123,  12'd59,  12'd50,  -12'd350,  -12'd394,  -12'd459,  12'd15,  12'd160,  12'd355,  12'd29,  -12'd137,  -12'd22,  -12'd58,  -12'd25,  -12'd50,  
12'd210,  -12'd303,  12'd248,  12'd15,  -12'd502,  12'd37,  -12'd727,  12'd103,  -12'd503,  12'd543,  -12'd56,  12'd187,  -12'd116,  -12'd98,  12'd170,  12'd353,  
-12'd203,  -12'd212,  -12'd171,  -12'd104,  12'd207,  -12'd166,  -12'd381,  -12'd102,  -12'd520,  -12'd91,  -12'd97,  -12'd68,  12'd110,  12'd131,  12'd269,  12'd205,  
-12'd65,  12'd155,  -12'd311,  -12'd36,  12'd113,  -12'd342,  -12'd157,  12'd107,  -12'd189,  -12'd308,  12'd18,  12'd217,  -12'd250,  -12'd266,  -12'd166,  -12'd19,  
-12'd922,  -12'd466,  12'd41,  -12'd157,  12'd268,  -12'd191,  -12'd320,  -12'd78,  12'd5,  12'd408,  -12'd183,  12'd162,  -12'd390,  -12'd156,  -12'd44,  -12'd441,  
-12'd574,  -12'd503,  -12'd87,  12'd430,  -12'd74,  -12'd103,  -12'd885,  12'd216,  12'd203,  12'd83,  12'd45,  -12'd191,  12'd39,  -12'd185,  -12'd58,  -12'd274,  
-12'd425,  -12'd330,  12'd485,  -12'd237,  12'd184,  -12'd127,  -12'd376,  -12'd205,  -12'd176,  12'd361,  12'd238,  12'd88,  -12'd51,  -12'd139,  -12'd270,  -12'd79,  
12'd163,  -12'd299,  12'd140,  12'd44,  -12'd181,  12'd161,  12'd190,  12'd130,  12'd165,  12'd82,  12'd147,  12'd117,  -12'd61,  -12'd124,  12'd20,  -12'd62,  
-12'd115,  -12'd0,  -12'd183,  12'd365,  12'd157,  12'd352,  12'd84,  12'd314,  -12'd21,  -12'd232,  12'd271,  12'd276,  12'd185,  12'd229,  12'd434,  12'd390,  
-12'd125,  -12'd96,  -12'd14,  12'd227,  -12'd35,  12'd81,  12'd300,  12'd265,  12'd460,  12'd263,  -12'd57,  12'd26,  -12'd265,  12'd159,  12'd205,  12'd70,  
-12'd259,  12'd51,  -12'd377,  12'd257,  12'd43,  12'd275,  -12'd18,  12'd142,  12'd897,  12'd282,  12'd308,  12'd407,  -12'd101,  -12'd262,  12'd190,  12'd84,  
-12'd74,  -12'd26,  -12'd117,  12'd406,  12'd196,  12'd46,  12'd1,  12'd127,  12'd223,  12'd91,  12'd117,  12'd169,  12'd377,  -12'd1077,  12'd98,  12'd277,  
12'd280,  12'd220,  -12'd282,  -12'd134,  12'd205,  12'd124,  -12'd155,  12'd223,  12'd241,  12'd188,  12'd71,  12'd30,  12'd512,  -12'd334,  -12'd31,  -12'd19,  
12'd440,  12'd245,  -12'd126,  -12'd122,  12'd21,  12'd157,  12'd177,  12'd273,  12'd215,  -12'd37,  -12'd127,  -12'd205,  12'd290,  12'd63,  -12'd78,  12'd120,  
12'd365,  12'd516,  12'd11,  12'd182,  -12'd241,  12'd234,  -12'd170,  12'd28,  12'd211,  -12'd155,  -12'd168,  12'd54,  12'd247,  12'd232,  12'd127,  12'd83,  

-12'd130,  12'd59,  12'd125,  12'd197,  -12'd196,  -12'd32,  -12'd45,  12'd4,  -12'd116,  12'd238,  12'd218,  -12'd190,  12'd218,  -12'd65,  -12'd33,  12'd231,  
12'd63,  12'd53,  12'd207,  -12'd167,  -12'd41,  -12'd76,  -12'd419,  -12'd247,  12'd374,  -12'd27,  -12'd155,  -12'd166,  12'd106,  -12'd215,  12'd29,  -12'd99,  
-12'd60,  12'd92,  12'd202,  -12'd221,  -12'd33,  12'd125,  -12'd187,  12'd32,  12'd44,  12'd256,  12'd110,  -12'd119,  -12'd313,  12'd79,  -12'd0,  -12'd384,  
-12'd216,  -12'd239,  -12'd152,  12'd20,  12'd200,  -12'd60,  12'd48,  -12'd136,  12'd39,  -12'd8,  -12'd33,  12'd253,  12'd2,  -12'd170,  12'd64,  -12'd388,  
12'd157,  12'd80,  -12'd213,  -12'd46,  -12'd81,  12'd47,  -12'd408,  -12'd213,  12'd155,  -12'd187,  12'd256,  -12'd25,  12'd160,  -12'd40,  12'd149,  -12'd47,  
-12'd180,  12'd218,  12'd60,  12'd10,  12'd33,  -12'd322,  -12'd262,  12'd38,  -12'd124,  12'd124,  12'd291,  -12'd156,  12'd320,  12'd32,  -12'd166,  12'd190,  
12'd349,  -12'd305,  -12'd176,  -12'd159,  -12'd170,  -12'd84,  12'd115,  12'd247,  -12'd148,  -12'd25,  -12'd351,  -12'd279,  -12'd127,  12'd163,  -12'd75,  -12'd80,  
12'd145,  -12'd132,  -12'd53,  -12'd235,  -12'd298,  -12'd103,  12'd74,  12'd109,  -12'd403,  12'd28,  -12'd312,  -12'd315,  12'd64,  -12'd191,  -12'd256,  -12'd281,  
-12'd69,  12'd78,  -12'd196,  12'd14,  -12'd458,  12'd79,  12'd92,  -12'd44,  -12'd109,  -12'd215,  12'd210,  -12'd262,  12'd23,  -12'd22,  12'd98,  12'd51,  
-12'd105,  12'd270,  -12'd249,  12'd130,  -12'd237,  -12'd110,  -12'd211,  -12'd153,  -12'd400,  -12'd8,  12'd329,  12'd156,  12'd43,  12'd19,  -12'd408,  12'd98,  
12'd97,  -12'd146,  -12'd393,  -12'd345,  12'd20,  -12'd45,  -12'd196,  -12'd247,  12'd14,  12'd121,  -12'd86,  12'd5,  -12'd340,  -12'd340,  12'd24,  12'd196,  
-12'd358,  -12'd301,  12'd255,  12'd23,  -12'd108,  -12'd294,  12'd296,  -12'd151,  12'd149,  -12'd52,  12'd260,  12'd58,  12'd164,  12'd25,  -12'd277,  -12'd321,  
-12'd102,  12'd83,  12'd36,  -12'd21,  12'd150,  12'd258,  -12'd229,  -12'd140,  -12'd232,  12'd288,  12'd43,  12'd70,  12'd38,  -12'd62,  -12'd161,  -12'd103,  
-12'd153,  -12'd60,  12'd70,  -12'd240,  -12'd158,  12'd244,  -12'd379,  12'd212,  -12'd337,  -12'd66,  12'd55,  12'd86,  12'd116,  -12'd68,  -12'd124,  -12'd14,  
-12'd66,  -12'd330,  -12'd84,  12'd45,  12'd183,  12'd201,  -12'd347,  -12'd191,  12'd150,  12'd239,  -12'd130,  -12'd19,  -12'd296,  12'd70,  12'd161,  -12'd183,  
-12'd155,  -12'd5,  12'd175,  12'd164,  12'd146,  12'd228,  12'd69,  -12'd310,  -12'd181,  -12'd151,  -12'd311,  -12'd141,  12'd104,  -12'd255,  -12'd242,  12'd318,  
12'd195,  12'd319,  12'd107,  -12'd36,  -12'd190,  -12'd90,  -12'd106,  -12'd124,  -12'd290,  -12'd162,  -12'd43,  -12'd280,  -12'd128,  12'd69,  12'd307,  12'd96,  
-12'd167,  12'd115,  -12'd23,  -12'd263,  -12'd297,  12'd175,  12'd44,  -12'd35,  12'd108,  -12'd79,  12'd14,  12'd102,  -12'd130,  12'd115,  -12'd66,  -12'd1,  
12'd131,  -12'd145,  -12'd234,  12'd103,  12'd12,  -12'd13,  -12'd88,  12'd106,  12'd349,  -12'd42,  12'd129,  -12'd164,  -12'd25,  12'd133,  -12'd7,  -12'd145,  
-12'd50,  -12'd313,  -12'd73,  -12'd95,  12'd114,  12'd112,  -12'd156,  12'd118,  -12'd50,  12'd148,  -12'd176,  12'd170,  12'd76,  -12'd179,  12'd104,  -12'd202,  
12'd7,  12'd132,  12'd389,  -12'd377,  12'd75,  -12'd132,  12'd279,  12'd22,  12'd249,  12'd121,  -12'd120,  12'd88,  12'd372,  -12'd199,  -12'd49,  -12'd75,  
-12'd205,  -12'd16,  -12'd36,  12'd128,  12'd184,  -12'd359,  12'd172,  -12'd270,  -12'd296,  12'd238,  -12'd204,  -12'd12,  12'd131,  -12'd21,  12'd24,  -12'd32,  
-12'd288,  12'd75,  -12'd59,  -12'd308,  12'd186,  -12'd307,  12'd16,  12'd255,  -12'd149,  -12'd16,  -12'd65,  12'd200,  12'd110,  -12'd7,  -12'd179,  12'd13,  
12'd83,  12'd57,  -12'd250,  12'd269,  12'd152,  -12'd153,  -12'd357,  -12'd46,  12'd306,  12'd292,  -12'd158,  12'd121,  -12'd221,  -12'd148,  12'd211,  12'd235,  
-12'd335,  12'd84,  -12'd77,  12'd166,  -12'd12,  12'd77,  12'd220,  12'd340,  -12'd11,  -12'd199,  12'd210,  12'd154,  12'd119,  12'd62,  -12'd107,  12'd177,  

12'd6,  12'd18,  -12'd405,  12'd82,  12'd169,  -12'd29,  12'd257,  12'd279,  12'd98,  -12'd326,  12'd405,  12'd143,  12'd503,  12'd98,  12'd259,  12'd443,  
12'd18,  12'd299,  -12'd439,  12'd226,  12'd65,  12'd233,  12'd77,  12'd220,  12'd273,  12'd95,  12'd350,  -12'd103,  12'd210,  -12'd452,  12'd313,  12'd144,  
-12'd531,  -12'd109,  12'd108,  -12'd152,  12'd237,  12'd134,  -12'd647,  -12'd18,  -12'd339,  -12'd447,  -12'd369,  -12'd102,  12'd371,  12'd234,  12'd67,  12'd324,  
-12'd9,  -12'd342,  -12'd208,  -12'd251,  -12'd262,  -12'd164,  12'd79,  12'd88,  -12'd138,  12'd185,  12'd131,  12'd142,  -12'd370,  -12'd179,  -12'd192,  -12'd641,  
-12'd2,  -12'd271,  -12'd52,  -12'd378,  -12'd424,  12'd40,  -12'd104,  -12'd21,  -12'd5,  -12'd55,  -12'd223,  -12'd8,  -12'd375,  12'd329,  -12'd507,  -12'd214,  
-12'd279,  12'd273,  12'd48,  -12'd62,  12'd142,  12'd162,  12'd480,  -12'd117,  12'd45,  -12'd36,  12'd367,  12'd63,  -12'd308,  -12'd132,  -12'd363,  -12'd246,  
12'd58,  -12'd35,  -12'd35,  12'd0,  12'd206,  12'd132,  12'd1,  12'd2,  12'd214,  12'd280,  12'd205,  -12'd141,  -12'd28,  -12'd131,  12'd267,  -12'd215,  
12'd20,  12'd22,  12'd36,  -12'd74,  12'd264,  -12'd208,  -12'd314,  12'd74,  -12'd281,  -12'd27,  -12'd26,  12'd110,  -12'd179,  12'd207,  12'd3,  12'd80,  
-12'd22,  -12'd317,  -12'd432,  -12'd179,  -12'd132,  -12'd449,  -12'd156,  -12'd402,  12'd253,  -12'd282,  -12'd308,  -12'd247,  -12'd546,  12'd251,  -12'd167,  -12'd173,  
-12'd474,  12'd119,  12'd185,  -12'd176,  -12'd194,  -12'd115,  -12'd193,  -12'd512,  -12'd492,  12'd169,  -12'd238,  12'd55,  -12'd564,  12'd532,  -12'd201,  -12'd108,  
-12'd85,  -12'd47,  -12'd365,  -12'd73,  12'd73,  12'd22,  12'd365,  -12'd385,  12'd57,  -12'd236,  -12'd162,  -12'd373,  -12'd1,  12'd35,  -12'd204,  12'd59,  
-12'd142,  12'd243,  -12'd91,  -12'd20,  12'd96,  -12'd0,  -12'd107,  12'd7,  12'd535,  12'd185,  -12'd227,  -12'd39,  12'd148,  -12'd79,  12'd268,  12'd268,  
-12'd22,  12'd164,  12'd12,  -12'd9,  -12'd131,  12'd145,  -12'd64,  -12'd30,  12'd443,  12'd225,  12'd249,  -12'd138,  12'd173,  12'd192,  -12'd197,  -12'd64,  
-12'd577,  12'd211,  -12'd606,  12'd530,  12'd9,  12'd222,  12'd214,  -12'd76,  12'd496,  -12'd296,  12'd730,  12'd119,  -12'd75,  12'd68,  -12'd172,  12'd240,  
-12'd524,  -12'd37,  12'd411,  12'd412,  -12'd63,  -12'd75,  -12'd31,  12'd149,  -12'd101,  -12'd67,  12'd815,  12'd39,  12'd479,  -12'd121,  12'd13,  12'd220,  
12'd555,  12'd108,  12'd286,  -12'd243,  -12'd351,  12'd308,  -12'd197,  -12'd57,  12'd31,  12'd36,  -12'd536,  -12'd259,  -12'd349,  12'd420,  12'd120,  -12'd470,  
12'd200,  -12'd50,  -12'd13,  -12'd96,  -12'd21,  -12'd369,  -12'd222,  -12'd144,  -12'd114,  -12'd36,  -12'd181,  -12'd98,  12'd93,  12'd233,  12'd519,  12'd335,  
12'd151,  -12'd303,  12'd109,  -12'd375,  12'd249,  12'd21,  12'd244,  -12'd344,  12'd64,  12'd350,  12'd336,  12'd36,  -12'd88,  -12'd95,  -12'd151,  12'd99,  
-12'd6,  12'd738,  -12'd231,  12'd172,  12'd112,  -12'd76,  12'd19,  12'd46,  12'd169,  -12'd298,  12'd399,  -12'd43,  12'd187,  12'd56,  12'd202,  12'd294,  
-12'd55,  -12'd205,  -12'd210,  12'd11,  12'd17,  -12'd373,  -12'd19,  -12'd229,  -12'd338,  12'd242,  12'd407,  -12'd332,  -12'd20,  12'd24,  12'd67,  12'd551,  
12'd87,  12'd161,  12'd383,  12'd352,  -12'd255,  12'd164,  -12'd402,  12'd237,  -12'd465,  -12'd44,  -12'd408,  -12'd334,  -12'd263,  12'd312,  12'd70,  -12'd488,  
12'd223,  -12'd135,  -12'd211,  -12'd117,  -12'd211,  12'd7,  -12'd28,  -12'd53,  -12'd315,  -12'd136,  12'd4,  -12'd333,  12'd105,  12'd317,  12'd212,  12'd47,  
12'd130,  -12'd88,  -12'd80,  12'd162,  12'd521,  -12'd202,  12'd369,  12'd315,  -12'd352,  -12'd439,  -12'd66,  -12'd331,  -12'd238,  -12'd183,  -12'd326,  12'd24,  
-12'd579,  12'd319,  12'd60,  -12'd66,  12'd28,  12'd135,  -12'd226,  12'd343,  -12'd60,  12'd233,  -12'd298,  -12'd498,  -12'd292,  12'd307,  -12'd448,  12'd13,  
-12'd576,  -12'd93,  12'd29,  12'd420,  12'd149,  -12'd66,  -12'd171,  -12'd57,  -12'd423,  12'd702,  12'd52,  -12'd122,  -12'd102,  -12'd58,  -12'd29,  12'd113,  

-12'd304,  -12'd114,  -12'd135,  -12'd64,  12'd274,  -12'd96,  12'd126,  12'd236,  -12'd89,  12'd6,  12'd333,  -12'd419,  -12'd14,  -12'd352,  12'd312,  12'd48,  
-12'd310,  -12'd92,  -12'd2,  12'd100,  12'd132,  -12'd76,  -12'd690,  -12'd11,  -12'd375,  12'd334,  -12'd491,  -12'd184,  12'd248,  -12'd627,  -12'd10,  12'd7,  
-12'd97,  -12'd378,  12'd278,  12'd448,  -12'd222,  12'd107,  12'd290,  12'd342,  -12'd159,  12'd315,  12'd310,  -12'd153,  -12'd277,  -12'd468,  12'd103,  12'd355,  
12'd394,  -12'd617,  -12'd233,  12'd192,  -12'd21,  12'd397,  12'd354,  12'd220,  12'd255,  -12'd151,  12'd73,  12'd191,  12'd311,  12'd541,  -12'd138,  -12'd192,  
-12'd428,  -12'd14,  12'd141,  -12'd259,  12'd133,  12'd212,  12'd68,  -12'd187,  12'd402,  -12'd273,  12'd160,  12'd161,  -12'd537,  12'd214,  -12'd45,  -12'd130,  
-12'd424,  12'd25,  -12'd341,  -12'd159,  -12'd208,  -12'd420,  -12'd502,  -12'd22,  -12'd126,  -12'd321,  12'd358,  -12'd16,  -12'd130,  -12'd213,  -12'd6,  12'd164,  
-12'd173,  -12'd260,  -12'd426,  -12'd392,  12'd270,  12'd59,  -12'd96,  12'd98,  -12'd98,  -12'd46,  12'd314,  12'd25,  -12'd169,  -12'd279,  12'd146,  12'd131,  
12'd224,  -12'd142,  -12'd278,  12'd140,  -12'd1,  -12'd112,  -12'd25,  -12'd20,  -12'd331,  12'd268,  -12'd29,  -12'd3,  -12'd102,  -12'd428,  12'd294,  12'd273,  
12'd520,  12'd48,  -12'd158,  -12'd40,  -12'd71,  -12'd232,  12'd359,  12'd227,  -12'd111,  12'd132,  -12'd100,  12'd38,  -12'd180,  12'd62,  12'd67,  12'd81,  
-12'd150,  12'd233,  -12'd82,  12'd272,  -12'd218,  12'd266,  12'd135,  -12'd99,  -12'd373,  -12'd10,  12'd47,  -12'd240,  12'd107,  12'd86,  -12'd168,  -12'd231,  
-12'd326,  -12'd108,  12'd62,  -12'd133,  -12'd367,  -12'd239,  12'd298,  12'd211,  12'd338,  -12'd191,  12'd260,  -12'd139,  -12'd307,  -12'd95,  12'd79,  -12'd326,  
12'd258,  -12'd240,  12'd117,  -12'd236,  -12'd468,  -12'd375,  12'd114,  -12'd103,  -12'd70,  12'd180,  -12'd338,  -12'd275,  12'd62,  12'd291,  12'd394,  -12'd270,  
12'd222,  -12'd113,  12'd298,  -12'd193,  -12'd323,  12'd75,  12'd55,  12'd76,  12'd70,  12'd67,  12'd22,  12'd187,  -12'd103,  12'd61,  -12'd156,  -12'd137,  
-12'd170,  -12'd36,  -12'd54,  12'd169,  12'd87,  12'd145,  12'd103,  12'd235,  12'd129,  12'd221,  12'd43,  12'd284,  -12'd79,  -12'd153,  12'd18,  12'd224,  
-12'd148,  -12'd14,  12'd92,  12'd78,  -12'd95,  -12'd126,  12'd121,  -12'd50,  12'd68,  12'd297,  12'd93,  -12'd195,  -12'd17,  -12'd64,  -12'd52,  -12'd217,  
-12'd346,  -12'd337,  12'd204,  12'd425,  -12'd22,  12'd303,  -12'd216,  12'd245,  12'd192,  12'd90,  12'd199,  -12'd90,  -12'd189,  12'd37,  12'd66,  12'd111,  
-12'd495,  -12'd139,  -12'd96,  12'd84,  12'd1,  -12'd212,  12'd229,  -12'd323,  -12'd205,  12'd431,  12'd313,  -12'd159,  -12'd213,  -12'd35,  12'd320,  -12'd107,  
-12'd52,  12'd211,  12'd107,  12'd135,  -12'd29,  12'd144,  12'd76,  12'd132,  -12'd122,  -12'd251,  -12'd263,  -12'd25,  -12'd6,  12'd89,  -12'd61,  -12'd270,  
12'd1,  -12'd46,  12'd313,  12'd366,  -12'd421,  -12'd141,  -12'd8,  -12'd162,  -12'd388,  -12'd245,  -12'd80,  12'd88,  12'd134,  -12'd14,  12'd37,  12'd323,  
12'd9,  12'd84,  12'd74,  12'd106,  -12'd186,  -12'd96,  12'd216,  12'd26,  -12'd234,  -12'd58,  12'd313,  -12'd161,  -12'd271,  12'd164,  -12'd337,  12'd176,  
-12'd202,  12'd175,  -12'd166,  12'd318,  -12'd147,  -12'd52,  12'd153,  12'd26,  12'd254,  12'd78,  12'd211,  -12'd122,  12'd161,  -12'd421,  -12'd98,  -12'd61,  
12'd78,  12'd264,  12'd165,  -12'd89,  12'd13,  12'd140,  -12'd95,  -12'd375,  12'd207,  12'd210,  12'd89,  12'd273,  12'd91,  -12'd321,  -12'd19,  12'd78,  
12'd14,  12'd118,  12'd111,  12'd224,  -12'd130,  12'd57,  12'd21,  -12'd63,  12'd449,  12'd31,  12'd126,  -12'd334,  12'd221,  -12'd9,  12'd297,  12'd44,  
12'd377,  -12'd76,  -12'd131,  -12'd2,  -12'd112,  12'd50,  12'd298,  -12'd15,  -12'd145,  -12'd96,  12'd388,  -12'd149,  12'd223,  12'd269,  -12'd326,  -12'd254,  
12'd135,  12'd141,  -12'd268,  -12'd16,  12'd63,  -12'd34,  -12'd129,  -12'd9,  12'd157,  -12'd131,  12'd130,  -12'd23,  -12'd245,  -12'd21,  -12'd73,  -12'd177,  

-12'd130,  12'd434,  12'd343,  12'd104,  -12'd102,  12'd155,  12'd157,  -12'd446,  12'd202,  -12'd297,  -12'd440,  12'd190,  -12'd193,  12'd192,  -12'd171,  -12'd137,  
-12'd45,  -12'd27,  12'd536,  -12'd486,  12'd57,  -12'd109,  -12'd49,  -12'd9,  12'd93,  -12'd90,  12'd95,  -12'd188,  12'd30,  12'd583,  12'd22,  -12'd235,  
-12'd473,  12'd108,  12'd175,  -12'd34,  -12'd182,  12'd99,  -12'd119,  12'd17,  12'd36,  -12'd232,  12'd172,  12'd120,  -12'd414,  12'd586,  -12'd76,  -12'd390,  
12'd89,  12'd5,  -12'd251,  12'd144,  -12'd65,  12'd299,  12'd120,  -12'd81,  12'd131,  12'd184,  -12'd352,  12'd119,  -12'd236,  12'd188,  -12'd250,  -12'd29,  
12'd287,  12'd147,  -12'd59,  12'd219,  -12'd121,  12'd61,  12'd244,  12'd12,  12'd336,  -12'd171,  -12'd39,  12'd181,  12'd292,  12'd284,  12'd21,  12'd260,  
12'd44,  12'd346,  12'd46,  12'd79,  -12'd311,  -12'd152,  12'd215,  12'd271,  -12'd191,  12'd466,  -12'd149,  12'd142,  -12'd172,  12'd466,  12'd280,  12'd120,  
12'd167,  12'd25,  12'd453,  -12'd281,  -12'd153,  -12'd397,  -12'd298,  12'd132,  12'd286,  -12'd39,  -12'd68,  -12'd193,  12'd267,  12'd530,  12'd275,  12'd296,  
12'd34,  -12'd311,  12'd327,  -12'd12,  -12'd13,  -12'd22,  -12'd278,  12'd144,  12'd259,  12'd49,  12'd175,  -12'd169,  -12'd112,  12'd38,  -12'd335,  -12'd317,  
-12'd201,  12'd173,  12'd265,  -12'd120,  12'd62,  12'd284,  -12'd136,  12'd50,  -12'd32,  12'd206,  -12'd231,  12'd207,  -12'd165,  -12'd91,  12'd72,  12'd107,  
12'd290,  -12'd275,  -12'd201,  12'd24,  -12'd95,  12'd166,  -12'd80,  -12'd314,  12'd149,  -12'd507,  -12'd127,  -12'd116,  -12'd321,  12'd96,  -12'd138,  12'd182,  
12'd407,  -12'd65,  -12'd9,  12'd414,  -12'd175,  12'd622,  -12'd405,  12'd186,  12'd154,  12'd38,  12'd260,  -12'd114,  12'd599,  12'd199,  -12'd62,  12'd173,  
-12'd110,  12'd354,  12'd60,  12'd173,  -12'd270,  12'd335,  -12'd72,  12'd432,  12'd147,  12'd281,  -12'd49,  -12'd61,  12'd127,  -12'd174,  12'd50,  -12'd364,  
12'd153,  -12'd40,  -12'd14,  12'd271,  -12'd70,  12'd406,  12'd150,  12'd138,  -12'd33,  -12'd104,  12'd425,  12'd15,  12'd389,  -12'd419,  -12'd210,  12'd11,  
-12'd28,  12'd68,  -12'd237,  12'd48,  12'd20,  -12'd233,  -12'd129,  -12'd230,  -12'd3,  -12'd290,  12'd396,  12'd210,  12'd15,  -12'd67,  12'd67,  -12'd78,  
-12'd123,  -12'd270,  -12'd45,  -12'd96,  -12'd109,  12'd24,  12'd181,  12'd157,  -12'd198,  -12'd235,  -12'd205,  -12'd18,  12'd543,  -12'd64,  -12'd64,  12'd459,  
12'd116,  12'd395,  -12'd168,  12'd9,  12'd742,  12'd150,  -12'd134,  -12'd189,  -12'd146,  12'd138,  -12'd58,  12'd426,  12'd206,  -12'd56,  12'd77,  12'd393,  
-12'd365,  -12'd53,  -12'd72,  -12'd12,  12'd175,  -12'd478,  12'd142,  12'd126,  -12'd74,  12'd80,  12'd82,  12'd81,  12'd105,  -12'd286,  -12'd143,  12'd101,  
-12'd56,  -12'd255,  12'd180,  12'd128,  12'd244,  -12'd145,  12'd144,  -12'd331,  12'd201,  12'd26,  -12'd104,  12'd80,  -12'd43,  12'd103,  -12'd276,  12'd26,  
12'd330,  12'd98,  12'd215,  12'd181,  -12'd163,  -12'd132,  12'd125,  -12'd29,  12'd260,  12'd371,  12'd300,  -12'd117,  -12'd32,  12'd312,  12'd24,  12'd363,  
-12'd180,  12'd204,  12'd127,  -12'd147,  -12'd241,  -12'd259,  -12'd379,  -12'd194,  -12'd389,  -12'd3,  -12'd98,  -12'd152,  -12'd249,  -12'd257,  12'd197,  12'd306,  
12'd147,  12'd364,  -12'd91,  -12'd232,  12'd236,  12'd125,  12'd77,  -12'd144,  12'd296,  -12'd334,  -12'd226,  12'd437,  -12'd315,  -12'd126,  -12'd134,  -12'd151,  
12'd85,  -12'd339,  -12'd61,  -12'd233,  12'd11,  -12'd122,  12'd421,  -12'd264,  -12'd30,  -12'd133,  -12'd83,  12'd33,  -12'd308,  -12'd115,  12'd301,  -12'd209,  
12'd327,  -12'd19,  12'd127,  -12'd123,  12'd159,  -12'd297,  12'd27,  -12'd114,  12'd36,  12'd131,  -12'd267,  -12'd242,  -12'd300,  12'd340,  -12'd78,  -12'd66,  
-12'd108,  12'd4,  -12'd26,  -12'd27,  -12'd181,  12'd28,  -12'd197,  12'd173,  12'd153,  12'd7,  -12'd22,  -12'd0,  -12'd204,  12'd474,  12'd304,  -12'd43,  
12'd64,  -12'd252,  12'd581,  12'd329,  12'd47,  12'd29,  12'd160,  12'd223,  -12'd91,  -12'd230,  -12'd214,  12'd77,  12'd297,  -12'd133,  12'd600,  12'd339,  

12'd151,  -12'd3,  -12'd248,  -12'd428,  -12'd418,  12'd382,  12'd310,  12'd73,  12'd400,  -12'd273,  12'd96,  12'd98,  -12'd66,  12'd231,  -12'd233,  -12'd21,  
-12'd48,  -12'd386,  -12'd240,  12'd116,  -12'd33,  12'd187,  -12'd237,  -12'd355,  -12'd62,  -12'd286,  12'd96,  -12'd9,  -12'd44,  -12'd137,  12'd300,  12'd177,  
12'd222,  12'd52,  -12'd175,  12'd184,  -12'd272,  12'd200,  -12'd123,  12'd110,  12'd82,  -12'd78,  12'd60,  -12'd257,  -12'd118,  -12'd293,  -12'd73,  -12'd12,  
-12'd299,  -12'd1,  -12'd34,  12'd286,  12'd204,  12'd132,  -12'd180,  -12'd227,  -12'd97,  12'd62,  12'd198,  -12'd112,  12'd215,  -12'd738,  12'd102,  12'd185,  
-12'd450,  -12'd446,  12'd143,  12'd62,  12'd252,  -12'd301,  -12'd158,  12'd156,  -12'd89,  -12'd252,  12'd176,  -12'd145,  12'd195,  12'd270,  -12'd94,  12'd483,  
12'd104,  12'd178,  -12'd66,  12'd277,  -12'd17,  12'd146,  -12'd341,  -12'd139,  -12'd346,  12'd491,  -12'd398,  12'd3,  -12'd161,  -12'd135,  12'd9,  12'd126,  
12'd144,  -12'd56,  12'd97,  12'd404,  -12'd336,  -12'd12,  -12'd577,  12'd252,  12'd270,  -12'd183,  -12'd81,  -12'd338,  12'd370,  12'd31,  12'd244,  12'd155,  
-12'd332,  12'd41,  12'd8,  -12'd198,  -12'd179,  12'd32,  12'd90,  12'd25,  12'd401,  12'd433,  12'd672,  -12'd139,  12'd67,  -12'd40,  -12'd137,  -12'd7,  
-12'd704,  -12'd328,  -12'd75,  -12'd193,  -12'd211,  -12'd129,  12'd203,  12'd238,  12'd73,  12'd508,  12'd12,  -12'd58,  12'd69,  -12'd135,  12'd263,  12'd100,  
-12'd248,  12'd2,  12'd103,  -12'd107,  -12'd284,  12'd132,  -12'd179,  -12'd62,  12'd216,  12'd148,  12'd264,  12'd182,  12'd155,  -12'd419,  12'd55,  12'd171,  
12'd214,  12'd4,  -12'd215,  -12'd41,  12'd247,  -12'd92,  -12'd801,  -12'd1,  12'd241,  12'd282,  12'd178,  -12'd138,  12'd192,  -12'd26,  -12'd55,  -12'd8,  
-12'd160,  12'd280,  12'd156,  -12'd265,  12'd17,  12'd116,  -12'd238,  12'd429,  12'd207,  12'd83,  -12'd211,  12'd218,  -12'd32,  12'd69,  -12'd53,  -12'd199,  
12'd201,  -12'd173,  -12'd305,  12'd109,  12'd345,  12'd122,  12'd58,  -12'd274,  -12'd25,  -12'd154,  12'd133,  12'd160,  12'd326,  -12'd185,  12'd175,  -12'd289,  
-12'd166,  12'd297,  12'd45,  -12'd164,  12'd122,  -12'd286,  -12'd42,  12'd132,  -12'd179,  12'd159,  12'd308,  -12'd53,  -12'd170,  -12'd42,  -12'd60,  -12'd100,  
12'd189,  12'd209,  -12'd106,  -12'd115,  12'd74,  12'd319,  12'd192,  12'd95,  12'd46,  -12'd7,  12'd127,  -12'd170,  12'd358,  -12'd136,  12'd120,  -12'd70,  
12'd160,  -12'd11,  12'd64,  12'd237,  12'd433,  12'd68,  12'd420,  -12'd200,  12'd478,  12'd307,  -12'd14,  -12'd111,  12'd106,  12'd228,  12'd181,  12'd365,  
12'd399,  12'd205,  12'd72,  12'd55,  -12'd111,  12'd66,  -12'd178,  -12'd84,  12'd103,  12'd182,  12'd186,  12'd457,  12'd501,  12'd50,  12'd97,  12'd238,  
-12'd82,  -12'd1,  -12'd42,  12'd284,  12'd86,  -12'd226,  12'd44,  -12'd227,  12'd116,  12'd377,  -12'd101,  -12'd221,  -12'd0,  -12'd307,  -12'd156,  12'd114,  
-12'd113,  -12'd102,  -12'd235,  -12'd143,  12'd126,  -12'd208,  12'd28,  -12'd173,  -12'd41,  12'd1,  -12'd261,  -12'd168,  -12'd255,  -12'd173,  12'd213,  12'd269,  
12'd240,  -12'd337,  12'd364,  12'd174,  -12'd90,  12'd358,  12'd10,  -12'd111,  12'd140,  12'd688,  12'd62,  -12'd293,  12'd65,  12'd273,  -12'd54,  12'd97,  
12'd38,  -12'd59,  -12'd68,  12'd263,  12'd137,  12'd181,  12'd293,  12'd403,  12'd308,  12'd245,  12'd192,  -12'd246,  12'd329,  -12'd112,  -12'd14,  -12'd123,  
12'd222,  -12'd483,  -12'd184,  -12'd246,  12'd235,  -12'd190,  -12'd134,  12'd55,  -12'd113,  -12'd82,  12'd24,  -12'd90,  12'd127,  12'd190,  -12'd24,  12'd54,  
-12'd308,  -12'd212,  -12'd216,  -12'd70,  12'd37,  12'd25,  -12'd167,  -12'd249,  12'd49,  12'd49,  -12'd126,  12'd424,  -12'd111,  12'd39,  12'd61,  -12'd44,  
12'd121,  -12'd68,  -12'd255,  12'd96,  12'd142,  -12'd85,  -12'd156,  -12'd14,  12'd209,  -12'd222,  12'd55,  -12'd166,  -12'd131,  12'd176,  -12'd155,  12'd232,  
-12'd13,  12'd42,  12'd55,  12'd193,  -12'd1,  12'd181,  -12'd18,  12'd204,  -12'd79,  -12'd121,  12'd212,  -12'd37,  12'd48,  -12'd154,  12'd210,  12'd357,  

-12'd222,  12'd121,  12'd244,  -12'd255,  12'd241,  -12'd410,  12'd96,  -12'd462,  12'd163,  12'd132,  12'd156,  -12'd226,  12'd132,  12'd461,  12'd97,  12'd290,  
-12'd344,  -12'd327,  12'd260,  -12'd21,  12'd33,  -12'd120,  12'd333,  -12'd354,  12'd24,  -12'd269,  12'd113,  12'd88,  -12'd183,  12'd481,  -12'd107,  12'd162,  
12'd276,  -12'd157,  12'd304,  -12'd223,  -12'd578,  12'd32,  -12'd26,  -12'd123,  -12'd239,  -12'd157,  12'd352,  -12'd392,  -12'd290,  12'd615,  12'd144,  -12'd203,  
12'd229,  12'd143,  -12'd245,  -12'd356,  -12'd168,  -12'd62,  12'd266,  12'd253,  12'd148,  -12'd68,  -12'd123,  12'd16,  12'd304,  -12'd304,  12'd230,  -12'd37,  
12'd130,  12'd852,  -12'd480,  12'd307,  -12'd93,  12'd105,  12'd183,  -12'd32,  -12'd37,  12'd12,  12'd426,  12'd88,  12'd579,  12'd124,  12'd18,  12'd529,  
-12'd303,  -12'd93,  12'd188,  -12'd132,  -12'd309,  -12'd257,  12'd266,  -12'd153,  -12'd201,  -12'd90,  12'd376,  -12'd15,  12'd105,  12'd271,  12'd115,  12'd134,  
12'd172,  12'd12,  -12'd95,  12'd144,  12'd239,  -12'd255,  12'd402,  12'd170,  -12'd5,  -12'd19,  12'd396,  12'd115,  12'd15,  12'd196,  -12'd334,  -12'd306,  
12'd58,  -12'd364,  12'd135,  -12'd410,  12'd63,  12'd36,  -12'd124,  12'd17,  12'd519,  -12'd14,  12'd75,  12'd64,  -12'd40,  -12'd153,  -12'd320,  -12'd186,  
12'd206,  12'd502,  12'd24,  12'd141,  12'd54,  -12'd4,  -12'd198,  12'd607,  12'd159,  12'd137,  12'd395,  -12'd62,  -12'd77,  -12'd145,  12'd93,  -12'd283,  
12'd43,  12'd98,  12'd127,  -12'd8,  12'd215,  12'd294,  -12'd29,  12'd356,  -12'd17,  12'd608,  12'd107,  12'd47,  -12'd78,  12'd207,  12'd455,  12'd4,  
12'd322,  12'd27,  12'd164,  -12'd174,  -12'd714,  12'd312,  12'd526,  -12'd137,  -12'd338,  12'd151,  12'd165,  12'd192,  -12'd80,  -12'd40,  12'd173,  12'd422,  
-12'd121,  12'd173,  12'd238,  12'd36,  12'd157,  -12'd166,  12'd102,  12'd125,  12'd2,  12'd18,  -12'd204,  -12'd85,  -12'd92,  12'd413,  -12'd47,  -12'd78,  
-12'd231,  12'd98,  12'd19,  -12'd239,  12'd176,  -12'd221,  -12'd141,  -12'd86,  -12'd122,  -12'd140,  -12'd2,  -12'd50,  12'd228,  -12'd85,  -12'd252,  12'd105,  
-12'd195,  -12'd183,  -12'd386,  -12'd81,  12'd98,  -12'd152,  -12'd434,  -12'd276,  -12'd179,  12'd355,  -12'd188,  12'd79,  -12'd88,  -12'd374,  12'd244,  12'd326,  
-12'd97,  12'd41,  12'd187,  -12'd5,  12'd233,  -12'd77,  -12'd327,  -12'd171,  12'd123,  12'd63,  12'd143,  12'd153,  -12'd22,  -12'd140,  12'd471,  12'd196,  
12'd42,  12'd111,  12'd414,  12'd44,  -12'd180,  12'd113,  -12'd55,  12'd562,  12'd52,  12'd15,  12'd97,  -12'd1,  -12'd13,  12'd20,  12'd191,  12'd64,  
-12'd124,  12'd189,  12'd101,  12'd410,  -12'd263,  12'd93,  -12'd30,  12'd3,  -12'd448,  -12'd213,  -12'd102,  -12'd349,  -12'd312,  12'd85,  12'd114,  -12'd380,  
12'd153,  -12'd271,  12'd161,  12'd137,  12'd288,  -12'd180,  12'd1,  12'd86,  12'd215,  -12'd297,  -12'd13,  -12'd49,  12'd264,  12'd258,  -12'd175,  -12'd323,  
12'd42,  -12'd72,  -12'd321,  -12'd91,  12'd395,  12'd286,  12'd34,  -12'd42,  12'd62,  12'd1,  12'd351,  12'd122,  12'd3,  12'd5,  -12'd30,  12'd13,  
12'd271,  12'd480,  12'd432,  -12'd275,  12'd87,  12'd62,  12'd187,  12'd36,  12'd73,  -12'd117,  -12'd16,  12'd255,  12'd89,  -12'd133,  12'd128,  -12'd2,  
-12'd429,  -12'd37,  -12'd39,  -12'd53,  -12'd114,  12'd223,  -12'd86,  12'd44,  12'd33,  -12'd19,  -12'd149,  12'd194,  -12'd227,  12'd117,  -12'd171,  12'd39,  
-12'd418,  -12'd153,  12'd90,  12'd259,  12'd194,  12'd430,  12'd366,  12'd20,  12'd266,  -12'd63,  12'd202,  -12'd66,  12'd347,  -12'd132,  -12'd59,  12'd22,  
-12'd247,  12'd55,  -12'd134,  12'd50,  12'd67,  12'd266,  12'd100,  12'd97,  12'd364,  -12'd94,  12'd395,  12'd60,  -12'd84,  -12'd168,  -12'd211,  12'd240,  
12'd471,  12'd51,  12'd438,  12'd88,  -12'd24,  -12'd128,  -12'd299,  12'd308,  -12'd39,  12'd125,  12'd242,  12'd245,  12'd141,  12'd79,  -12'd454,  -12'd219,  
12'd348,  12'd19,  12'd258,  -12'd36,  12'd170,  -12'd68,  12'd189,  -12'd118,  12'd388,  12'd171,  -12'd155,  12'd574,  12'd187,  -12'd344,  12'd2,  -12'd63,  

-12'd407,  -12'd54,  -12'd208,  12'd39,  12'd133,  12'd42,  -12'd336,  12'd314,  -12'd210,  12'd69,  -12'd67,  -12'd350,  12'd547,  -12'd74,  -12'd65,  -12'd356,  
-12'd126,  12'd186,  12'd31,  -12'd13,  12'd199,  12'd229,  -12'd189,  12'd9,  12'd127,  12'd112,  -12'd340,  -12'd65,  12'd181,  -12'd68,  12'd208,  12'd41,  
-12'd267,  -12'd70,  12'd429,  12'd56,  -12'd349,  12'd178,  12'd168,  -12'd292,  12'd24,  -12'd196,  12'd68,  -12'd196,  -12'd147,  12'd336,  12'd247,  12'd398,  
-12'd93,  -12'd187,  12'd22,  12'd454,  -12'd397,  -12'd290,  -12'd202,  -12'd5,  12'd447,  12'd109,  12'd272,  12'd10,  -12'd274,  12'd42,  12'd58,  -12'd117,  
-12'd9,  -12'd280,  12'd195,  -12'd135,  12'd366,  -12'd262,  -12'd219,  -12'd237,  -12'd79,  -12'd142,  12'd281,  12'd53,  -12'd87,  12'd53,  -12'd41,  12'd30,  
-12'd332,  -12'd101,  -12'd478,  12'd277,  12'd189,  -12'd389,  -12'd87,  -12'd399,  12'd60,  -12'd268,  12'd251,  -12'd117,  12'd120,  -12'd17,  -12'd319,  12'd154,  
-12'd219,  -12'd245,  -12'd421,  12'd239,  12'd496,  -12'd207,  -12'd201,  -12'd86,  -12'd142,  12'd186,  -12'd200,  12'd286,  12'd339,  -12'd199,  -12'd12,  12'd229,  
-12'd54,  12'd71,  12'd47,  12'd147,  12'd94,  -12'd103,  -12'd6,  -12'd38,  -12'd167,  12'd6,  12'd187,  12'd130,  12'd246,  -12'd56,  -12'd490,  -12'd25,  
-12'd25,  12'd30,  12'd105,  -12'd215,  -12'd114,  12'd243,  -12'd206,  -12'd200,  -12'd183,  12'd185,  12'd215,  12'd42,  12'd114,  12'd442,  -12'd11,  -12'd39,  
12'd139,  12'd427,  12'd333,  12'd219,  -12'd97,  -12'd271,  12'd254,  -12'd23,  12'd213,  12'd199,  12'd53,  12'd4,  -12'd252,  12'd261,  12'd440,  -12'd143,  
-12'd197,  12'd133,  -12'd308,  -12'd355,  -12'd229,  12'd286,  -12'd462,  12'd127,  12'd360,  -12'd217,  12'd403,  12'd113,  -12'd46,  -12'd20,  12'd217,  12'd217,  
12'd220,  12'd44,  12'd7,  12'd89,  12'd108,  12'd212,  -12'd183,  -12'd322,  12'd112,  12'd560,  12'd51,  12'd56,  12'd135,  -12'd335,  -12'd299,  12'd475,  
12'd159,  12'd136,  -12'd391,  12'd130,  12'd462,  -12'd354,  12'd41,  12'd156,  -12'd168,  12'd166,  12'd324,  12'd306,  12'd33,  -12'd129,  12'd4,  12'd398,  
12'd67,  12'd193,  12'd186,  12'd87,  12'd199,  -12'd117,  12'd183,  12'd164,  12'd293,  12'd299,  12'd285,  -12'd133,  -12'd235,  12'd41,  -12'd342,  -12'd438,  
12'd251,  12'd109,  12'd43,  12'd208,  -12'd396,  12'd244,  12'd86,  -12'd69,  12'd114,  -12'd255,  -12'd299,  -12'd42,  12'd319,  -12'd223,  -12'd504,  -12'd45,  
12'd18,  -12'd80,  -12'd246,  -12'd40,  -12'd375,  -12'd134,  -12'd262,  -12'd132,  12'd165,  -12'd16,  12'd375,  -12'd122,  -12'd78,  -12'd304,  12'd30,  12'd185,  
-12'd231,  12'd11,  -12'd331,  12'd159,  12'd137,  -12'd12,  -12'd242,  12'd372,  -12'd124,  12'd64,  12'd200,  12'd253,  12'd116,  -12'd174,  12'd107,  12'd252,  
12'd180,  12'd311,  -12'd366,  12'd106,  12'd182,  12'd75,  -12'd68,  12'd69,  12'd81,  -12'd234,  12'd203,  12'd263,  12'd147,  12'd209,  -12'd154,  -12'd68,  
12'd98,  -12'd110,  -12'd344,  12'd440,  12'd73,  -12'd198,  -12'd45,  12'd22,  12'd98,  -12'd203,  12'd394,  -12'd149,  12'd251,  -12'd7,  12'd53,  12'd233,  
12'd207,  -12'd172,  -12'd314,  12'd169,  12'd340,  12'd302,  -12'd60,  -12'd179,  12'd240,  -12'd33,  12'd38,  12'd21,  12'd615,  12'd62,  -12'd29,  12'd60,  
-12'd39,  -12'd170,  -12'd86,  -12'd254,  -12'd73,  -12'd8,  12'd374,  -12'd362,  -12'd342,  12'd266,  12'd142,  -12'd147,  12'd219,  12'd9,  12'd180,  12'd215,  
-12'd25,  12'd383,  12'd143,  -12'd109,  12'd30,  -12'd456,  -12'd77,  -12'd1,  -12'd9,  -12'd128,  12'd342,  -12'd161,  12'd1,  -12'd513,  12'd56,  12'd146,  
12'd210,  12'd140,  -12'd184,  -12'd18,  12'd258,  -12'd85,  -12'd127,  -12'd170,  -12'd205,  12'd514,  -12'd182,  -12'd13,  12'd174,  -12'd95,  12'd192,  -12'd235,  
-12'd312,  12'd452,  -12'd43,  12'd162,  12'd15,  -12'd248,  -12'd119,  -12'd25,  -12'd25,  12'd38,  12'd28,  -12'd405,  12'd378,  12'd63,  -12'd130,  -12'd252,  
12'd47,  12'd335,  12'd114,  -12'd157,  -12'd57,  12'd225,  -12'd465,  12'd213,  12'd99,  12'd332,  -12'd336,  12'd125,  -12'd160,  -12'd163,  12'd59,  -12'd108,  

12'd107,  12'd1,  -12'd240,  -12'd27,  -12'd32,  12'd58,  12'd3,  -12'd116,  12'd259,  -12'd115,  -12'd150,  12'd138,  12'd204,  -12'd63,  -12'd279,  12'd158,  
12'd279,  -12'd110,  12'd125,  12'd158,  -12'd272,  12'd126,  -12'd31,  12'd23,  -12'd375,  12'd172,  -12'd301,  -12'd8,  -12'd302,  -12'd250,  -12'd343,  -12'd183,  
-12'd114,  -12'd235,  -12'd74,  -12'd24,  12'd32,  12'd40,  -12'd8,  -12'd187,  12'd128,  -12'd173,  -12'd54,  -12'd228,  -12'd139,  -12'd126,  -12'd138,  12'd126,  
-12'd213,  -12'd141,  -12'd182,  12'd0,  -12'd15,  -12'd52,  12'd65,  12'd123,  12'd98,  -12'd180,  -12'd71,  12'd154,  -12'd136,  -12'd328,  -12'd31,  -12'd141,  
12'd32,  12'd168,  12'd189,  -12'd185,  -12'd53,  -12'd185,  -12'd58,  12'd3,  12'd105,  12'd7,  -12'd299,  -12'd13,  12'd24,  12'd122,  12'd272,  12'd152,  
-12'd119,  -12'd131,  -12'd118,  -12'd162,  12'd39,  12'd134,  -12'd234,  -12'd211,  12'd6,  -12'd360,  12'd179,  12'd32,  -12'd177,  12'd176,  -12'd100,  -12'd92,  
12'd243,  12'd2,  12'd149,  -12'd195,  12'd166,  -12'd245,  -12'd17,  -12'd170,  -12'd136,  -12'd157,  12'd132,  12'd11,  12'd251,  -12'd69,  12'd78,  12'd135,  
12'd35,  -12'd217,  -12'd171,  -12'd96,  12'd120,  -12'd50,  -12'd423,  12'd203,  -12'd91,  12'd9,  12'd87,  -12'd327,  12'd252,  -12'd52,  -12'd57,  -12'd265,  
12'd300,  -12'd112,  12'd11,  -12'd10,  12'd42,  12'd331,  -12'd277,  12'd112,  -12'd243,  -12'd187,  -12'd96,  12'd74,  12'd217,  -12'd161,  12'd220,  12'd132,  
12'd257,  -12'd52,  12'd140,  12'd363,  -12'd35,  -12'd165,  -12'd356,  12'd291,  12'd40,  -12'd368,  -12'd93,  -12'd37,  -12'd53,  -12'd22,  12'd233,  12'd231,  
-12'd27,  12'd32,  -12'd67,  -12'd136,  -12'd360,  12'd73,  -12'd191,  -12'd91,  -12'd178,  -12'd382,  -12'd78,  12'd17,  12'd56,  -12'd42,  12'd201,  -12'd335,  
12'd249,  -12'd90,  12'd245,  12'd164,  -12'd425,  12'd178,  -12'd78,  12'd92,  -12'd358,  12'd328,  12'd173,  12'd18,  12'd155,  -12'd191,  12'd21,  12'd44,  
12'd3,  -12'd171,  -12'd281,  -12'd24,  12'd12,  -12'd369,  12'd60,  -12'd79,  12'd171,  12'd75,  -12'd129,  12'd91,  -12'd63,  12'd44,  12'd154,  12'd126,  
-12'd116,  12'd129,  -12'd189,  -12'd3,  -12'd14,  -12'd179,  -12'd164,  -12'd219,  -12'd367,  -12'd364,  -12'd177,  -12'd195,  -12'd204,  12'd59,  -12'd169,  -12'd67,  
-12'd238,  12'd17,  -12'd270,  -12'd186,  -12'd150,  -12'd54,  -12'd19,  -12'd347,  -12'd16,  -12'd161,  -12'd316,  -12'd80,  12'd7,  -12'd38,  12'd147,  12'd17,  
-12'd100,  -12'd6,  -12'd37,  -12'd25,  12'd79,  -12'd141,  -12'd130,  12'd43,  12'd219,  -12'd125,  -12'd177,  -12'd110,  -12'd158,  -12'd65,  12'd156,  12'd247,  
12'd167,  12'd307,  12'd135,  -12'd215,  -12'd45,  12'd237,  -12'd379,  -12'd10,  12'd65,  -12'd90,  12'd81,  12'd34,  -12'd22,  12'd102,  -12'd191,  12'd171,  
-12'd364,  12'd15,  -12'd38,  12'd39,  -12'd269,  12'd250,  12'd146,  -12'd6,  -12'd298,  -12'd217,  -12'd0,  -12'd140,  -12'd264,  -12'd123,  12'd90,  -12'd30,  
12'd265,  -12'd25,  -12'd167,  12'd188,  12'd265,  12'd145,  -12'd26,  -12'd182,  12'd236,  -12'd97,  -12'd145,  12'd30,  12'd337,  12'd62,  12'd103,  -12'd17,  
12'd299,  -12'd322,  -12'd132,  -12'd192,  -12'd96,  -12'd115,  -12'd171,  -12'd21,  -12'd206,  12'd177,  12'd44,  12'd37,  -12'd78,  12'd275,  -12'd138,  12'd178,  
-12'd74,  12'd124,  -12'd6,  12'd288,  -12'd371,  12'd153,  12'd95,  -12'd77,  12'd33,  -12'd300,  -12'd37,  -12'd243,  12'd141,  -12'd275,  -12'd300,  -12'd368,  
-12'd104,  12'd23,  -12'd158,  12'd298,  12'd93,  -12'd383,  -12'd56,  -12'd171,  12'd96,  12'd190,  12'd110,  12'd122,  -12'd422,  -12'd111,  -12'd135,  -12'd250,  
-12'd71,  12'd12,  -12'd302,  -12'd161,  12'd55,  12'd74,  -12'd196,  -12'd183,  12'd31,  -12'd302,  12'd286,  -12'd359,  -12'd119,  -12'd306,  12'd202,  -12'd266,  
-12'd186,  -12'd121,  12'd67,  -12'd88,  -12'd191,  12'd353,  -12'd26,  -12'd117,  -12'd65,  12'd228,  -12'd179,  12'd163,  -12'd232,  -12'd86,  12'd75,  -12'd215,  
12'd48,  12'd84,  12'd13,  -12'd57,  12'd88,  -12'd205,  12'd2,  -12'd227,  12'd322,  -12'd193,  12'd257,  -12'd174,  -12'd322,  -12'd39,  12'd27,  -12'd127,  

-12'd221,  -12'd32,  -12'd154,  -12'd5,  12'd90,  12'd216,  12'd83,  -12'd237,  -12'd409,  12'd1,  -12'd75,  12'd211,  -12'd124,  -12'd206,  -12'd266,  -12'd178,  
12'd28,  -12'd84,  -12'd369,  -12'd22,  -12'd124,  12'd75,  -12'd71,  12'd105,  -12'd16,  12'd77,  12'd96,  12'd185,  -12'd253,  -12'd499,  -12'd111,  12'd79,  
-12'd428,  -12'd207,  -12'd130,  -12'd97,  12'd521,  12'd131,  -12'd200,  -12'd246,  -12'd318,  12'd160,  12'd70,  -12'd20,  12'd411,  -12'd808,  -12'd66,  -12'd6,  
-12'd487,  -12'd417,  12'd163,  12'd118,  12'd28,  -12'd397,  -12'd36,  12'd65,  -12'd252,  -12'd5,  -12'd106,  12'd185,  12'd59,  -12'd9,  12'd94,  -12'd140,  
-12'd92,  -12'd116,  -12'd43,  -12'd222,  12'd358,  -12'd144,  -12'd162,  12'd273,  12'd178,  -12'd147,  12'd69,  12'd144,  -12'd155,  -12'd94,  -12'd97,  -12'd41,  
-12'd367,  12'd153,  12'd21,  -12'd211,  -12'd270,  -12'd356,  -12'd1,  12'd188,  12'd347,  -12'd160,  12'd478,  12'd167,  12'd119,  12'd108,  12'd53,  12'd67,  
12'd45,  12'd243,  12'd205,  12'd34,  12'd43,  -12'd307,  12'd148,  -12'd243,  -12'd13,  12'd294,  -12'd357,  12'd211,  12'd224,  -12'd215,  12'd359,  12'd217,  
-12'd212,  -12'd220,  -12'd362,  -12'd7,  12'd169,  -12'd135,  12'd38,  -12'd191,  -12'd97,  -12'd88,  12'd49,  12'd321,  12'd266,  -12'd550,  12'd279,  -12'd6,  
12'd126,  -12'd92,  -12'd103,  12'd88,  -12'd85,  -12'd39,  12'd206,  12'd194,  12'd241,  12'd35,  12'd42,  12'd125,  12'd277,  12'd247,  12'd148,  12'd392,  
12'd231,  12'd169,  12'd102,  12'd428,  12'd23,  12'd184,  12'd42,  12'd132,  -12'd178,  -12'd460,  -12'd22,  -12'd11,  12'd80,  12'd153,  -12'd169,  -12'd6,  
12'd58,  12'd25,  -12'd222,  -12'd90,  12'd135,  -12'd57,  -12'd486,  12'd24,  12'd181,  12'd142,  -12'd382,  -12'd173,  12'd368,  12'd187,  12'd167,  12'd134,  
-12'd11,  12'd148,  -12'd218,  12'd65,  -12'd43,  -12'd208,  -12'd367,  -12'd82,  -12'd299,  12'd117,  12'd320,  -12'd293,  -12'd25,  12'd222,  12'd161,  -12'd17,  
12'd272,  -12'd343,  12'd102,  12'd293,  -12'd221,  12'd147,  -12'd251,  -12'd14,  -12'd304,  12'd115,  12'd126,  12'd385,  -12'd59,  -12'd626,  12'd19,  -12'd111,  
12'd206,  -12'd459,  -12'd94,  -12'd37,  12'd347,  -12'd183,  12'd144,  -12'd202,  12'd10,  12'd337,  -12'd170,  12'd90,  12'd165,  12'd49,  12'd46,  12'd242,  
-12'd145,  -12'd212,  -12'd91,  -12'd268,  12'd285,  -12'd46,  12'd231,  -12'd471,  -12'd172,  12'd150,  12'd145,  -12'd268,  -12'd19,  -12'd14,  12'd59,  12'd463,  
-12'd406,  -12'd131,  -12'd402,  -12'd146,  12'd265,  -12'd364,  -12'd316,  -12'd166,  -12'd53,  -12'd40,  -12'd147,  -12'd111,  -12'd227,  -12'd231,  -12'd203,  12'd136,  
12'd305,  12'd134,  -12'd74,  12'd318,  12'd522,  -12'd204,  -12'd273,  -12'd297,  12'd313,  12'd182,  -12'd245,  12'd36,  12'd34,  -12'd464,  -12'd126,  12'd73,  
-12'd96,  12'd191,  12'd192,  12'd203,  -12'd308,  12'd229,  -12'd102,  12'd259,  12'd59,  -12'd94,  12'd79,  -12'd51,  -12'd138,  -12'd653,  12'd256,  -12'd60,  
12'd94,  12'd235,  -12'd109,  -12'd79,  -12'd46,  -12'd94,  12'd130,  12'd114,  12'd425,  -12'd173,  -12'd14,  12'd137,  12'd115,  12'd281,  -12'd116,  -12'd126,  
-12'd27,  12'd42,  -12'd96,  -12'd70,  -12'd427,  -12'd229,  12'd266,  -12'd436,  12'd283,  -12'd130,  12'd132,  -12'd415,  -12'd228,  -12'd181,  -12'd248,  -12'd184,  
12'd120,  -12'd52,  -12'd171,  -12'd361,  -12'd176,  -12'd51,  12'd198,  -12'd178,  12'd477,  -12'd22,  12'd387,  12'd223,  12'd248,  -12'd391,  12'd179,  12'd26,  
12'd419,  -12'd259,  -12'd98,  -12'd18,  12'd120,  12'd60,  -12'd51,  12'd124,  12'd245,  12'd189,  12'd108,  12'd246,  -12'd100,  -12'd50,  -12'd249,  -12'd28,  
12'd77,  12'd188,  12'd272,  -12'd21,  -12'd384,  -12'd29,  12'd223,  12'd272,  12'd387,  12'd446,  12'd134,  12'd195,  12'd292,  12'd180,  12'd48,  -12'd109,  
12'd98,  -12'd127,  12'd200,  -12'd61,  -12'd194,  -12'd191,  12'd116,  -12'd35,  -12'd133,  -12'd228,  12'd62,  12'd242,  12'd116,  12'd400,  -12'd264,  12'd255,  
-12'd16,  -12'd237,  12'd230,  -12'd128,  -12'd322,  12'd46,  12'd77,  -12'd33,  12'd337,  -12'd111,  12'd1,  -12'd85,  -12'd38,  12'd127,  -12'd53,  -12'd187,  

12'd247,  -12'd235,  -12'd59,  -12'd418,  -12'd79,  -12'd74,  -12'd299,  12'd5,  12'd208,  12'd258,  -12'd21,  -12'd93,  -12'd22,  12'd3,  12'd107,  12'd34,  
12'd307,  -12'd68,  12'd92,  -12'd159,  12'd257,  12'd42,  -12'd173,  -12'd221,  12'd199,  -12'd422,  -12'd101,  -12'd315,  -12'd330,  -12'd69,  -12'd73,  12'd177,  
-12'd241,  -12'd119,  -12'd52,  12'd295,  -12'd132,  12'd179,  12'd283,  12'd310,  -12'd417,  -12'd287,  -12'd172,  -12'd177,  -12'd295,  12'd173,  12'd28,  12'd103,  
12'd64,  12'd210,  12'd113,  -12'd118,  12'd97,  -12'd27,  12'd286,  -12'd135,  -12'd147,  12'd37,  12'd131,  -12'd72,  12'd308,  -12'd143,  12'd47,  -12'd132,  
-12'd66,  12'd230,  12'd95,  -12'd247,  -12'd267,  12'd270,  -12'd74,  -12'd26,  -12'd188,  12'd88,  12'd30,  -12'd294,  12'd44,  -12'd25,  -12'd280,  12'd216,  
-12'd102,  12'd4,  -12'd150,  -12'd99,  -12'd165,  -12'd268,  -12'd268,  -12'd81,  12'd124,  -12'd239,  -12'd264,  -12'd9,  12'd297,  -12'd157,  -12'd204,  -12'd195,  
12'd97,  -12'd177,  12'd354,  12'd288,  -12'd112,  -12'd48,  -12'd201,  -12'd324,  12'd246,  -12'd0,  -12'd147,  12'd65,  12'd10,  12'd27,  -12'd325,  -12'd423,  
-12'd69,  12'd161,  12'd88,  12'd47,  12'd130,  -12'd72,  -12'd180,  -12'd109,  -12'd287,  -12'd53,  -12'd45,  12'd196,  12'd284,  12'd90,  -12'd202,  -12'd110,  
12'd184,  -12'd159,  -12'd109,  -12'd179,  12'd350,  12'd275,  -12'd176,  -12'd278,  -12'd192,  -12'd347,  12'd175,  -12'd178,  12'd24,  12'd85,  -12'd181,  -12'd73,  
-12'd200,  -12'd191,  12'd234,  -12'd241,  12'd199,  -12'd74,  12'd261,  -12'd242,  12'd93,  -12'd24,  -12'd54,  -12'd168,  -12'd309,  12'd130,  -12'd230,  12'd145,  
-12'd230,  -12'd254,  12'd85,  12'd147,  12'd28,  -12'd57,  -12'd82,  -12'd91,  -12'd45,  -12'd227,  -12'd446,  -12'd266,  12'd155,  12'd230,  12'd166,  -12'd39,  
12'd150,  12'd227,  -12'd164,  -12'd132,  -12'd92,  12'd11,  12'd208,  -12'd68,  -12'd59,  -12'd291,  12'd77,  12'd112,  12'd96,  -12'd197,  -12'd391,  12'd7,  
12'd57,  -12'd302,  12'd2,  -12'd158,  -12'd74,  -12'd174,  12'd112,  -12'd224,  12'd78,  12'd20,  -12'd10,  -12'd76,  -12'd235,  -12'd70,  -12'd75,  12'd304,  
-12'd184,  -12'd328,  12'd34,  -12'd22,  12'd130,  -12'd195,  -12'd42,  -12'd244,  -12'd374,  -12'd112,  -12'd204,  12'd50,  -12'd299,  -12'd65,  12'd7,  12'd94,  
-12'd116,  -12'd134,  -12'd17,  -12'd97,  12'd52,  12'd4,  12'd189,  12'd7,  12'd323,  -12'd11,  12'd116,  -12'd189,  -12'd9,  12'd82,  12'd318,  -12'd93,  
12'd108,  12'd207,  12'd188,  12'd152,  -12'd291,  12'd244,  12'd363,  -12'd132,  12'd255,  -12'd92,  -12'd132,  -12'd154,  12'd136,  -12'd359,  12'd6,  -12'd351,  
12'd119,  -12'd10,  -12'd217,  12'd68,  -12'd80,  -12'd182,  12'd35,  12'd275,  -12'd27,  12'd208,  12'd295,  -12'd326,  12'd192,  -12'd314,  12'd192,  12'd149,  
-12'd58,  -12'd281,  -12'd417,  12'd252,  12'd71,  -12'd121,  12'd161,  -12'd277,  12'd182,  12'd150,  -12'd80,  12'd53,  -12'd187,  12'd58,  -12'd110,  -12'd10,  
-12'd371,  -12'd104,  -12'd56,  12'd22,  12'd6,  -12'd151,  -12'd117,  12'd19,  -12'd68,  -12'd81,  12'd86,  12'd333,  -12'd271,  -12'd16,  12'd2,  12'd13,  
-12'd362,  12'd142,  12'd294,  -12'd199,  -12'd217,  12'd13,  -12'd271,  12'd220,  -12'd344,  12'd14,  12'd197,  -12'd55,  12'd77,  -12'd63,  12'd132,  -12'd170,  
-12'd26,  -12'd352,  -12'd253,  -12'd3,  -12'd104,  -12'd150,  -12'd214,  -12'd341,  12'd141,  -12'd58,  -12'd28,  -12'd135,  -12'd301,  12'd179,  -12'd111,  -12'd20,  
12'd105,  12'd274,  12'd49,  -12'd19,  12'd111,  -12'd38,  12'd49,  -12'd88,  12'd329,  -12'd5,  12'd182,  12'd127,  -12'd2,  12'd126,  12'd54,  -12'd0,  
12'd222,  -12'd103,  -12'd27,  -12'd385,  12'd71,  -12'd110,  12'd218,  -12'd112,  12'd10,  12'd104,  -12'd271,  -12'd138,  -12'd4,  12'd60,  -12'd89,  -12'd348,  
12'd78,  -12'd39,  12'd118,  -12'd152,  12'd14,  -12'd209,  12'd325,  -12'd187,  -12'd92,  -12'd4,  12'd84,  -12'd64,  -12'd233,  -12'd96,  -12'd174,  -12'd118,  
12'd276,  12'd73,  12'd122,  -12'd58,  -12'd156,  12'd137,  12'd191,  12'd50,  12'd55,  -12'd227,  12'd213,  -12'd91,  12'd63,  -12'd101,  -12'd247,  -12'd179,  

12'd59,  -12'd159,  12'd166,  -12'd149,  -12'd244,  -12'd40,  -12'd192,  -12'd62,  -12'd159,  12'd263,  12'd158,  -12'd7,  12'd198,  -12'd79,  -12'd192,  -12'd387,  
-12'd104,  12'd159,  -12'd231,  -12'd224,  -12'd300,  12'd187,  12'd164,  -12'd372,  12'd9,  -12'd223,  -12'd95,  -12'd149,  12'd24,  -12'd41,  12'd53,  12'd105,  
-12'd9,  12'd363,  12'd70,  -12'd110,  -12'd2,  12'd196,  12'd41,  -12'd204,  12'd271,  12'd303,  12'd4,  -12'd128,  -12'd325,  -12'd136,  -12'd203,  12'd22,  
12'd69,  -12'd317,  -12'd278,  12'd280,  12'd217,  12'd313,  12'd164,  -12'd265,  -12'd116,  12'd156,  -12'd294,  12'd126,  -12'd151,  -12'd376,  -12'd342,  -12'd131,  
12'd197,  -12'd60,  -12'd67,  -12'd233,  12'd287,  12'd91,  12'd31,  -12'd118,  12'd99,  12'd161,  -12'd58,  -12'd64,  -12'd322,  -12'd10,  12'd186,  12'd84,  
-12'd257,  12'd276,  -12'd349,  -12'd338,  -12'd460,  12'd18,  -12'd17,  -12'd317,  12'd153,  -12'd332,  -12'd321,  -12'd177,  -12'd198,  12'd87,  -12'd71,  -12'd70,  
-12'd257,  -12'd131,  -12'd251,  12'd201,  -12'd81,  -12'd363,  -12'd280,  -12'd153,  -12'd139,  -12'd463,  -12'd249,  -12'd259,  -12'd211,  -12'd137,  -12'd97,  -12'd232,  
-12'd164,  -12'd3,  -12'd330,  -12'd212,  -12'd96,  -12'd155,  12'd222,  -12'd176,  -12'd298,  12'd338,  -12'd203,  -12'd127,  12'd18,  -12'd437,  -12'd235,  12'd136,  
-12'd15,  -12'd202,  12'd44,  -12'd301,  -12'd268,  -12'd215,  -12'd12,  -12'd247,  12'd131,  -12'd73,  -12'd173,  12'd22,  12'd18,  -12'd224,  12'd28,  -12'd39,  
12'd2,  -12'd404,  12'd228,  -12'd152,  12'd183,  12'd148,  12'd256,  -12'd58,  12'd34,  12'd132,  -12'd157,  -12'd12,  12'd106,  -12'd63,  12'd237,  12'd42,  
-12'd338,  12'd158,  -12'd62,  -12'd292,  -12'd157,  -12'd208,  -12'd215,  12'd172,  12'd122,  12'd250,  -12'd163,  -12'd233,  -12'd45,  12'd68,  12'd258,  -12'd67,  
-12'd192,  -12'd125,  -12'd307,  -12'd56,  -12'd2,  12'd72,  -12'd128,  -12'd474,  12'd146,  -12'd107,  -12'd124,  12'd96,  -12'd136,  -12'd247,  12'd1,  -12'd48,  
12'd74,  -12'd338,  -12'd167,  12'd125,  12'd178,  12'd60,  12'd72,  -12'd66,  -12'd420,  -12'd173,  12'd77,  -12'd32,  -12'd153,  12'd57,  -12'd165,  12'd32,  
12'd65,  -12'd88,  -12'd471,  12'd10,  12'd100,  -12'd84,  12'd10,  12'd42,  -12'd39,  12'd88,  12'd71,  -12'd114,  -12'd156,  12'd258,  12'd35,  12'd49,  
-12'd111,  -12'd40,  -12'd84,  -12'd80,  12'd108,  -12'd156,  -12'd45,  -12'd235,  12'd15,  -12'd247,  -12'd334,  12'd167,  12'd217,  12'd123,  -12'd197,  12'd42,  
-12'd284,  12'd60,  -12'd7,  -12'd279,  12'd2,  -12'd82,  12'd11,  -12'd280,  -12'd119,  -12'd104,  -12'd28,  -12'd187,  -12'd105,  12'd73,  -12'd94,  12'd137,  
-12'd0,  -12'd7,  -12'd9,  -12'd80,  12'd19,  -12'd304,  -12'd26,  12'd56,  -12'd336,  12'd201,  12'd10,  -12'd333,  -12'd309,  12'd187,  12'd303,  12'd130,  
-12'd323,  -12'd155,  12'd106,  -12'd98,  -12'd71,  -12'd281,  -12'd88,  12'd231,  12'd396,  12'd130,  -12'd396,  -12'd217,  -12'd155,  12'd38,  12'd60,  -12'd156,  
-12'd201,  12'd236,  -12'd496,  -12'd168,  -12'd162,  -12'd58,  12'd22,  -12'd104,  -12'd309,  -12'd193,  -12'd340,  12'd98,  -12'd17,  -12'd121,  -12'd292,  -12'd52,  
12'd44,  -12'd333,  -12'd103,  -12'd284,  -12'd20,  -12'd157,  -12'd133,  -12'd304,  -12'd51,  -12'd74,  -12'd210,  -12'd350,  12'd50,  -12'd11,  12'd79,  12'd172,  
-12'd206,  -12'd8,  -12'd171,  -12'd455,  -12'd102,  -12'd84,  12'd89,  12'd102,  12'd104,  -12'd380,  -12'd56,  -12'd101,  12'd60,  -12'd8,  12'd42,  -12'd112,  
12'd212,  -12'd112,  -12'd214,  -12'd241,  -12'd138,  12'd178,  12'd140,  -12'd324,  12'd167,  12'd49,  12'd95,  12'd16,  12'd40,  12'd119,  12'd4,  -12'd247,  
12'd113,  -12'd113,  -12'd330,  12'd203,  12'd172,  12'd148,  12'd58,  -12'd207,  -12'd105,  12'd54,  12'd295,  12'd21,  -12'd20,  -12'd274,  12'd0,  12'd160,  
12'd192,  -12'd248,  -12'd159,  -12'd93,  -12'd163,  -12'd258,  -12'd169,  -12'd134,  12'd168,  -12'd251,  -12'd66,  -12'd2,  -12'd15,  12'd11,  12'd26,  12'd59,  
-12'd74,  12'd141,  -12'd72,  -12'd91,  12'd122,  -12'd178,  -12'd316,  -12'd205,  12'd45,  -12'd347,  12'd261,  -12'd146,  -12'd312,  -12'd146,  12'd99,  12'd128,  

12'd197,  12'd252,  12'd558,  12'd334,  -12'd47,  12'd24,  -12'd368,  12'd23,  -12'd94,  12'd206,  -12'd99,  -12'd36,  12'd241,  12'd182,  12'd322,  -12'd186,  
12'd265,  12'd156,  -12'd163,  -12'd10,  12'd367,  -12'd351,  12'd148,  -12'd145,  12'd571,  -12'd268,  -12'd42,  12'd416,  12'd108,  -12'd250,  -12'd251,  12'd46,  
12'd191,  12'd357,  -12'd270,  -12'd1,  -12'd198,  12'd374,  12'd81,  -12'd176,  -12'd276,  -12'd114,  -12'd184,  12'd5,  12'd65,  12'd456,  12'd50,  12'd190,  
12'd27,  12'd17,  12'd260,  -12'd15,  12'd67,  -12'd389,  -12'd52,  -12'd136,  12'd135,  -12'd49,  -12'd33,  12'd146,  12'd136,  12'd430,  -12'd217,  12'd187,  
12'd65,  12'd405,  -12'd422,  -12'd128,  12'd53,  -12'd58,  12'd268,  -12'd124,  12'd254,  12'd252,  12'd193,  12'd280,  -12'd101,  12'd424,  12'd77,  12'd7,  
-12'd194,  -12'd142,  12'd331,  -12'd42,  12'd79,  12'd23,  12'd254,  12'd338,  -12'd87,  12'd315,  12'd271,  -12'd65,  12'd144,  12'd157,  -12'd84,  12'd34,  
-12'd263,  -12'd135,  12'd252,  -12'd88,  -12'd290,  12'd68,  12'd191,  12'd75,  -12'd28,  12'd195,  12'd39,  -12'd55,  12'd155,  -12'd170,  12'd1,  -12'd358,  
12'd35,  12'd299,  -12'd19,  -12'd209,  12'd55,  -12'd217,  12'd148,  -12'd293,  12'd36,  -12'd0,  -12'd188,  12'd394,  12'd352,  -12'd79,  12'd33,  -12'd55,  
12'd211,  12'd182,  -12'd200,  12'd110,  12'd68,  -12'd13,  12'd68,  -12'd507,  12'd36,  -12'd525,  -12'd241,  12'd139,  -12'd21,  12'd264,  -12'd192,  12'd132,  
-12'd28,  12'd166,  -12'd512,  -12'd190,  12'd312,  -12'd176,  12'd202,  -12'd186,  12'd186,  -12'd85,  12'd203,  12'd199,  12'd313,  -12'd148,  12'd23,  -12'd98,  
12'd127,  12'd11,  12'd91,  12'd264,  -12'd267,  -12'd60,  12'd261,  12'd32,  -12'd8,  12'd208,  12'd181,  -12'd58,  12'd45,  12'd161,  12'd360,  12'd248,  
12'd108,  12'd6,  12'd110,  -12'd104,  -12'd30,  -12'd39,  12'd278,  12'd207,  12'd209,  12'd142,  12'd346,  -12'd125,  12'd41,  -12'd370,  12'd48,  -12'd110,  
12'd349,  -12'd379,  12'd215,  12'd461,  12'd200,  12'd256,  -12'd397,  12'd114,  12'd30,  12'd241,  12'd57,  12'd255,  12'd225,  12'd350,  12'd262,  12'd199,  
12'd299,  -12'd488,  -12'd255,  -12'd190,  12'd285,  -12'd97,  12'd166,  -12'd267,  -12'd199,  -12'd95,  -12'd258,  12'd164,  12'd283,  12'd103,  -12'd62,  -12'd215,  
12'd85,  -12'd319,  -12'd208,  12'd28,  -12'd149,  12'd1,  -12'd222,  -12'd303,  12'd2,  12'd264,  -12'd181,  12'd154,  -12'd121,  12'd262,  -12'd44,  12'd333,  
12'd118,  -12'd19,  12'd128,  -12'd177,  12'd298,  -12'd372,  12'd427,  -12'd26,  -12'd195,  12'd13,  12'd30,  12'd148,  12'd153,  12'd10,  -12'd16,  12'd287,  
12'd185,  -12'd251,  -12'd303,  -12'd1,  -12'd217,  12'd59,  12'd175,  12'd85,  12'd356,  12'd319,  -12'd224,  -12'd186,  -12'd126,  12'd324,  -12'd50,  12'd117,  
-12'd173,  12'd231,  -12'd139,  12'd175,  -12'd193,  12'd127,  12'd87,  -12'd63,  -12'd15,  -12'd220,  12'd293,  12'd247,  12'd98,  -12'd275,  -12'd148,  12'd34,  
-12'd43,  -12'd225,  -12'd102,  12'd121,  12'd425,  -12'd43,  -12'd25,  -12'd2,  -12'd62,  -12'd92,  12'd279,  -12'd186,  -12'd58,  -12'd92,  -12'd40,  -12'd265,  
-12'd85,  -12'd235,  -12'd235,  12'd161,  12'd467,  12'd41,  12'd102,  12'd77,  12'd104,  12'd327,  12'd7,  12'd277,  12'd74,  -12'd195,  -12'd102,  12'd306,  
12'd210,  12'd391,  -12'd120,  -12'd352,  -12'd59,  -12'd210,  -12'd6,  -12'd132,  -12'd445,  -12'd274,  12'd32,  -12'd15,  -12'd57,  12'd239,  12'd0,  -12'd275,  
-12'd169,  -12'd156,  12'd450,  12'd26,  -12'd108,  -12'd238,  -12'd330,  12'd197,  -12'd399,  -12'd360,  -12'd376,  -12'd147,  -12'd169,  12'd769,  -12'd151,  -12'd98,  
-12'd152,  12'd187,  12'd112,  -12'd56,  12'd85,  12'd0,  -12'd0,  -12'd42,  -12'd176,  -12'd257,  -12'd21,  -12'd111,  -12'd56,  12'd313,  12'd302,  -12'd280,  
-12'd269,  -12'd218,  -12'd304,  -12'd229,  -12'd204,  12'd367,  -12'd124,  12'd83,  -12'd129,  -12'd232,  12'd196,  12'd58,  12'd165,  12'd427,  12'd500,  12'd402,  
-12'd555,  12'd242,  12'd38,  12'd336,  -12'd76,  -12'd106,  12'd20,  -12'd33,  -12'd380,  -12'd53,  12'd279,  12'd157,  -12'd172,  -12'd51,  12'd494,  12'd157
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule



module bias_fc2_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC2-1][0:`OUTPUT_NUM_FC2-1][`WD_BIAS:0] weight	 = {
		24'd376858,  24'd432250,  24'd29999,  -24'd21180,  24'd203900,  -24'd35257,  24'd214653,  -24'd285062,  24'd149942,  24'd172424,  24'd241287,  24'd324760,  24'd306054,  24'd109385,  24'd386902,  24'd1789,  
24'd28800,  24'd347429,  24'd509845,  24'd403218,  24'd55283,  24'd293083,  -24'd21746,  -24'd254371,  -24'd400996,  -24'd132702,  -24'd107502,  -24'd140243,  -24'd206663,  -24'd140441,  24'd143746,  24'd39439,  
24'd236044,  24'd268803,  24'd150150,  24'd385287,  -24'd213047,  24'd26023,  -24'd343539,  24'd332436,  -24'd397889,  -24'd209506,  -24'd133163,  24'd243649,  -24'd9532,  24'd307082,  -24'd132963,  -24'd159572,  
-24'd53911,  24'd55608,  -24'd63297,  24'd287278,  24'd231376,  24'd227915,  -24'd149391,  24'd406123,  -24'd279679,  24'd37076,  24'd251134,  24'd110896,  -24'd132970,  24'd307661,  24'd327144,  24'd66815,  
24'd131364,  24'd119973,  -24'd302322,  24'd158931,  24'd47008,  -24'd154135,  -24'd42487,  24'd329397,  24'd366838,  24'd373655,  24'd391455,  24'd142308,  24'd61661,  24'd27682,  24'd173948,  -24'd11642,  
24'd233626,  -24'd79977,  24'd87200,  24'd305044
	 };
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule


module wieght_fc2_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2*`OUTPUT_BATCH_FC2)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC1*`OUTPUT_NUM_FC2 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC2*`KERNEL_SIZEX_FC2*`KERNEL_SIZEY_FC2-1][0:`OUTPUT_NUM_FC2-1][0:`OUTPUT_NUM_FC1-1][`WD:0] weight	 = {
12'd42,  -12'd168,  -12'd273,  12'd389,  12'd518,  -12'd105,  12'd217,  12'd408,  -12'd345,  -12'd64,  -12'd391,  12'd405,  -12'd279,  -12'd94,  12'd467,  12'd145,  
12'd217,  -12'd29,  -12'd19,  12'd233,  12'd255,  -12'd476,  12'd31,  12'd483,  12'd21,  -12'd49,  -12'd117,  -12'd46,  -12'd171,  12'd141,  12'd104,  -12'd214,  
12'd190,  12'd331,  -12'd259,  12'd149,  -12'd92,  12'd83,  12'd129,  12'd356,  -12'd89,  -12'd361,  12'd100,  12'd171,  12'd299,  12'd81,  -12'd430,  -12'd164,  
-12'd100,  12'd95,  12'd76,  12'd191,  -12'd188,  12'd134,  -12'd307,  12'd24,  12'd248,  -12'd256,  12'd16,  -12'd150,  12'd34,  12'd344,  -12'd86,  12'd232,  
12'd26,  12'd270,  12'd169,  -12'd199,  -12'd61,  -12'd225,  -12'd110,  12'd56,  12'd174,  12'd441,  -12'd218,  -12'd292,  12'd186,  -12'd92,  -12'd268,  12'd223,  
-12'd63,  -12'd39,  12'd111,  12'd16,  12'd158,  -12'd335,  -12'd247,  12'd64,  -12'd293,  12'd136,  -12'd348,  -12'd321,  12'd188,  12'd129,  12'd337,  -12'd165,  
-12'd24,  -12'd211,  -12'd74,  12'd609,  -12'd80,  -12'd238,  12'd30,  -12'd63,  -12'd290,  -12'd155,  -12'd380,  12'd426,  -12'd246,  -12'd238,  12'd109,  12'd217,  
12'd185,  12'd79,  -12'd299,  -12'd14,  12'd192,  -12'd39,  -12'd358,  -12'd235,  
-12'd180,  -12'd230,  12'd74,  12'd23,  -12'd36,  -12'd200,  -12'd362,  -12'd411,  12'd67,  12'd56,  12'd94,  -12'd449,  12'd4,  12'd74,  12'd341,  12'd207,  
-12'd13,  -12'd129,  12'd339,  -12'd147,  -12'd26,  12'd346,  12'd79,  -12'd166,  12'd75,  -12'd310,  -12'd101,  -12'd170,  12'd182,  12'd216,  12'd204,  12'd10,  
-12'd106,  -12'd41,  12'd423,  12'd181,  12'd101,  12'd67,  -12'd75,  -12'd24,  12'd276,  -12'd378,  12'd145,  12'd72,  12'd168,  -12'd10,  -12'd247,  -12'd395,  
12'd92,  -12'd359,  -12'd32,  12'd106,  12'd397,  12'd225,  -12'd346,  -12'd143,  -12'd158,  12'd236,  -12'd205,  12'd218,  12'd336,  12'd143,  12'd78,  12'd68,  
12'd124,  12'd35,  12'd88,  12'd12,  -12'd221,  12'd41,  -12'd252,  12'd17,  -12'd339,  -12'd200,  12'd38,  -12'd64,  -12'd181,  -12'd263,  12'd103,  -12'd133,  
12'd18,  -12'd36,  12'd314,  -12'd93,  -12'd17,  -12'd249,  -12'd17,  12'd11,  -12'd7,  -12'd36,  -12'd251,  12'd230,  12'd295,  12'd217,  -12'd283,  12'd103,  
12'd326,  12'd309,  -12'd189,  12'd45,  12'd188,  -12'd98,  12'd185,  -12'd557,  12'd273,  12'd44,  -12'd206,  -12'd373,  -12'd29,  12'd175,  -12'd347,  12'd301,  
12'd53,  -12'd22,  -12'd169,  -12'd10,  12'd251,  12'd72,  12'd352,  -12'd112,  
-12'd327,  -12'd161,  12'd164,  12'd237,  -12'd53,  12'd210,  12'd52,  12'd126,  -12'd235,  12'd7,  12'd18,  -12'd128,  12'd41,  12'd191,  -12'd17,  12'd191,  
-12'd240,  12'd98,  -12'd207,  12'd35,  12'd79,  12'd205,  -12'd64,  12'd119,  -12'd282,  -12'd269,  -12'd137,  12'd175,  -12'd58,  12'd109,  -12'd78,  12'd321,  
-12'd129,  12'd288,  12'd250,  12'd268,  -12'd268,  12'd343,  -12'd82,  12'd216,  12'd357,  12'd143,  -12'd137,  -12'd116,  -12'd96,  12'd401,  12'd74,  -12'd234,  
12'd33,  -12'd353,  12'd394,  12'd60,  12'd46,  -12'd491,  12'd304,  12'd131,  -12'd22,  12'd243,  12'd283,  12'd263,  12'd222,  -12'd120,  -12'd305,  -12'd71,  
-12'd200,  12'd39,  -12'd43,  -12'd142,  -12'd10,  -12'd169,  -12'd49,  12'd209,  -12'd63,  12'd160,  12'd261,  -12'd193,  -12'd349,  -12'd156,  12'd97,  -12'd291,  
12'd152,  -12'd315,  -12'd368,  -12'd92,  12'd221,  12'd99,  12'd267,  12'd141,  12'd20,  -12'd212,  12'd97,  -12'd185,  -12'd377,  12'd430,  12'd158,  -12'd12,  
-12'd287,  -12'd13,  12'd9,  -12'd20,  -12'd159,  12'd157,  -12'd279,  12'd298,  12'd28,  12'd222,  12'd124,  12'd93,  -12'd81,  -12'd12,  12'd264,  12'd140,  
12'd49,  12'd21,  12'd30,  -12'd50,  12'd480,  -12'd182,  -12'd15,  12'd169,  
12'd143,  -12'd37,  12'd91,  -12'd15,  12'd233,  12'd96,  12'd95,  -12'd247,  -12'd355,  12'd18,  -12'd370,  -12'd260,  12'd163,  12'd63,  12'd84,  12'd127,  
12'd329,  12'd152,  -12'd104,  -12'd304,  12'd152,  12'd171,  12'd285,  12'd46,  12'd197,  -12'd327,  12'd13,  -12'd537,  12'd109,  12'd3,  12'd273,  12'd515,  
12'd65,  12'd6,  12'd81,  12'd61,  12'd363,  -12'd135,  -12'd407,  12'd224,  -12'd144,  12'd96,  12'd175,  -12'd429,  12'd255,  12'd128,  -12'd547,  -12'd151,  
-12'd97,  12'd327,  12'd366,  12'd31,  -12'd94,  12'd57,  12'd19,  -12'd12,  12'd207,  12'd291,  -12'd10,  12'd9,  12'd115,  -12'd179,  12'd84,  -12'd330,  
-12'd103,  12'd49,  -12'd107,  12'd326,  -12'd408,  12'd30,  -12'd466,  -12'd8,  12'd203,  -12'd352,  -12'd45,  12'd186,  -12'd386,  -12'd138,  12'd296,  12'd94,  
-12'd121,  -12'd181,  12'd203,  -12'd65,  -12'd270,  12'd110,  12'd76,  -12'd243,  -12'd123,  -12'd98,  12'd269,  -12'd166,  12'd129,  -12'd13,  12'd318,  -12'd75,  
12'd273,  -12'd30,  12'd69,  -12'd133,  12'd330,  12'd454,  -12'd65,  -12'd855,  12'd58,  -12'd140,  -12'd184,  -12'd121,  12'd28,  -12'd557,  -12'd258,  12'd352,  
12'd24,  12'd23,  12'd35,  -12'd351,  -12'd397,  -12'd175,  12'd69,  12'd365,  
-12'd195,  -12'd37,  -12'd264,  -12'd151,  12'd187,  12'd249,  12'd191,  -12'd94,  -12'd90,  12'd198,  -12'd383,  12'd208,  12'd192,  12'd151,  12'd76,  12'd13,  
12'd144,  -12'd37,  12'd198,  -12'd207,  -12'd21,  12'd258,  12'd148,  12'd20,  12'd128,  -12'd307,  -12'd47,  12'd227,  12'd79,  -12'd128,  12'd184,  -12'd144,  
-12'd224,  12'd227,  -12'd120,  -12'd38,  -12'd34,  12'd9,  -12'd80,  12'd411,  -12'd410,  -12'd31,  -12'd592,  -12'd136,  12'd109,  12'd200,  12'd415,  12'd241,  
12'd222,  -12'd307,  -12'd333,  12'd325,  12'd47,  12'd298,  12'd122,  -12'd182,  -12'd94,  -12'd50,  12'd170,  -12'd101,  -12'd17,  12'd263,  12'd162,  -12'd165,  
12'd335,  -12'd136,  12'd186,  -12'd349,  12'd484,  -12'd84,  -12'd127,  12'd301,  12'd10,  -12'd1,  -12'd197,  -12'd3,  12'd80,  12'd34,  -12'd112,  12'd286,  
-12'd13,  -12'd191,  12'd294,  -12'd310,  -12'd102,  -12'd86,  -12'd74,  12'd38,  -12'd317,  12'd164,  12'd126,  12'd122,  12'd218,  -12'd262,  -12'd87,  -12'd63,  
-12'd116,  12'd69,  12'd158,  -12'd420,  -12'd11,  12'd1,  12'd221,  -12'd176,  -12'd66,  -12'd15,  -12'd165,  12'd692,  12'd189,  -12'd110,  -12'd368,  -12'd73,  
12'd385,  -12'd169,  12'd308,  -12'd196,  -12'd99,  12'd217,  12'd17,  -12'd194,  
-12'd361,  -12'd16,  12'd333,  12'd26,  -12'd402,  12'd405,  12'd139,  -12'd306,  -12'd72,  12'd203,  12'd550,  -12'd309,  -12'd194,  12'd2,  -12'd94,  -12'd37,  
-12'd38,  -12'd19,  -12'd184,  12'd148,  12'd84,  12'd224,  12'd296,  -12'd7,  -12'd28,  12'd50,  12'd226,  -12'd10,  -12'd166,  12'd291,  -12'd251,  -12'd42,  
-12'd204,  12'd97,  12'd48,  -12'd87,  12'd218,  12'd106,  -12'd238,  -12'd375,  12'd179,  12'd40,  -12'd118,  12'd351,  -12'd377,  12'd10,  -12'd74,  12'd112,  
12'd263,  12'd65,  12'd187,  12'd319,  12'd399,  12'd66,  12'd436,  12'd50,  -12'd529,  12'd76,  -12'd200,  -12'd53,  12'd320,  12'd50,  12'd231,  -12'd297,  
-12'd107,  -12'd300,  -12'd272,  12'd132,  -12'd379,  12'd242,  -12'd22,  -12'd27,  12'd68,  12'd278,  12'd111,  12'd156,  -12'd285,  12'd52,  -12'd97,  12'd155,  
12'd175,  -12'd95,  12'd77,  -12'd414,  12'd147,  12'd417,  12'd126,  -12'd214,  -12'd34,  12'd15,  12'd226,  12'd37,  -12'd29,  12'd164,  12'd91,  12'd210,  
12'd253,  12'd143,  12'd246,  -12'd97,  12'd232,  -12'd238,  12'd343,  12'd245,  12'd41,  -12'd167,  12'd48,  -12'd107,  -12'd247,  12'd3,  12'd305,  -12'd129,  
-12'd11,  12'd285,  12'd545,  12'd282,  -12'd106,  -12'd284,  -12'd219,  -12'd79,  
12'd121,  -12'd175,  12'd199,  -12'd154,  -12'd261,  -12'd340,  -12'd450,  12'd184,  -12'd468,  -12'd131,  -12'd333,  -12'd235,  -12'd167,  12'd207,  -12'd305,  12'd138,  
-12'd89,  12'd67,  12'd10,  -12'd94,  12'd177,  -12'd303,  -12'd46,  12'd185,  12'd206,  12'd227,  12'd204,  -12'd193,  -12'd67,  12'd47,  -12'd86,  12'd323,  
-12'd120,  12'd166,  12'd318,  12'd89,  12'd474,  -12'd129,  -12'd406,  -12'd335,  12'd1,  -12'd177,  -12'd76,  -12'd30,  -12'd319,  -12'd110,  -12'd272,  -12'd794,  
12'd83,  12'd74,  -12'd11,  12'd195,  12'd58,  12'd150,  12'd167,  12'd204,  12'd220,  12'd134,  12'd85,  12'd330,  12'd283,  -12'd599,  -12'd114,  12'd69,  
12'd62,  12'd68,  -12'd274,  -12'd203,  -12'd420,  12'd393,  -12'd50,  12'd60,  -12'd239,  12'd19,  12'd41,  -12'd190,  12'd204,  12'd206,  12'd138,  12'd55,  
-12'd120,  -12'd343,  -12'd32,  12'd171,  -12'd157,  -12'd300,  -12'd196,  -12'd91,  -12'd133,  12'd183,  12'd16,  -12'd203,  12'd133,  12'd289,  -12'd308,  12'd418,  
-12'd145,  -12'd224,  -12'd117,  -12'd141,  -12'd142,  12'd47,  12'd402,  12'd100,  -12'd260,  -12'd315,  -12'd10,  12'd164,  -12'd133,  -12'd178,  -12'd123,  12'd112,  
-12'd121,  12'd177,  -12'd404,  -12'd99,  12'd295,  12'd125,  12'd12,  -12'd110,  
12'd215,  -12'd63,  -12'd201,  -12'd237,  12'd239,  12'd131,  -12'd285,  -12'd71,  -12'd124,  -12'd131,  -12'd335,  12'd181,  12'd230,  -12'd45,  12'd357,  12'd52,  
12'd122,  12'd141,  -12'd118,  12'd21,  -12'd300,  12'd148,  -12'd119,  12'd478,  12'd115,  12'd417,  -12'd137,  -12'd313,  12'd367,  -12'd49,  12'd168,  12'd125,  
12'd155,  -12'd32,  -12'd98,  12'd47,  12'd347,  -12'd66,  12'd258,  -12'd25,  -12'd192,  -12'd144,  12'd28,  -12'd295,  12'd378,  12'd161,  -12'd69,  -12'd335,  
12'd62,  12'd171,  12'd168,  -12'd433,  -12'd45,  12'd120,  12'd364,  12'd89,  12'd21,  12'd211,  -12'd232,  12'd180,  12'd145,  12'd187,  12'd107,  -12'd168,  
12'd6,  12'd215,  12'd241,  -12'd76,  12'd101,  -12'd466,  12'd376,  12'd88,  12'd521,  -12'd328,  -12'd42,  -12'd477,  12'd111,  -12'd122,  12'd78,  12'd154,  
-12'd40,  -12'd278,  -12'd370,  12'd291,  -12'd151,  -12'd37,  12'd64,  -12'd47,  -12'd452,  -12'd314,  12'd343,  12'd61,  12'd404,  -12'd336,  -12'd37,  -12'd180,  
-12'd148,  12'd201,  -12'd175,  12'd357,  12'd94,  -12'd214,  -12'd293,  -12'd93,  -12'd199,  12'd125,  -12'd79,  12'd78,  -12'd244,  -12'd95,  -12'd35,  12'd279,  
-12'd261,  -12'd154,  -12'd11,  12'd217,  12'd138,  12'd291,  -12'd14,  12'd208,  
12'd65,  12'd169,  -12'd227,  -12'd38,  -12'd270,  12'd130,  -12'd362,  -12'd23,  -12'd163,  -12'd241,  -12'd177,  12'd242,  -12'd77,  12'd483,  -12'd46,  12'd50,  
12'd67,  -12'd472,  12'd229,  12'd302,  12'd109,  12'd329,  12'd13,  -12'd196,  12'd15,  -12'd236,  -12'd166,  12'd17,  -12'd123,  12'd141,  -12'd456,  -12'd77,  
-12'd40,  12'd172,  -12'd142,  -12'd98,  12'd23,  12'd190,  -12'd382,  12'd103,  -12'd237,  12'd140,  -12'd216,  -12'd156,  12'd157,  12'd273,  -12'd177,  12'd99,  
12'd82,  12'd182,  -12'd93,  12'd57,  12'd297,  12'd158,  -12'd263,  12'd26,  -12'd168,  12'd218,  12'd349,  12'd79,  -12'd390,  12'd204,  12'd364,  12'd338,  
12'd195,  -12'd210,  12'd97,  -12'd219,  12'd201,  12'd69,  12'd44,  -12'd265,  12'd265,  12'd283,  -12'd149,  12'd51,  -12'd165,  -12'd170,  12'd89,  -12'd106,  
12'd164,  -12'd253,  12'd122,  -12'd26,  -12'd252,  -12'd52,  -12'd161,  12'd47,  -12'd109,  -12'd160,  -12'd30,  12'd71,  12'd140,  -12'd67,  -12'd149,  -12'd269,  
12'd39,  -12'd75,  12'd497,  -12'd214,  12'd84,  -12'd388,  -12'd37,  -12'd107,  12'd234,  -12'd153,  -12'd395,  12'd78,  -12'd135,  -12'd51,  -12'd66,  12'd228,  
12'd244,  12'd168,  12'd230,  12'd125,  -12'd342,  -12'd143,  12'd161,  12'd411,  
-12'd253,  12'd37,  -12'd121,  12'd60,  12'd194,  12'd44,  12'd176,  12'd594,  -12'd195,  12'd103,  12'd244,  -12'd64,  -12'd90,  -12'd150,  12'd162,  -12'd88,  
-12'd77,  12'd251,  12'd196,  -12'd207,  12'd68,  -12'd142,  12'd192,  -12'd79,  12'd118,  12'd185,  -12'd40,  12'd117,  12'd37,  12'd326,  12'd143,  -12'd148,  
-12'd146,  12'd412,  -12'd217,  12'd135,  -12'd13,  -12'd645,  -12'd227,  12'd308,  -12'd483,  -12'd163,  12'd123,  12'd418,  12'd694,  12'd306,  -12'd32,  -12'd128,  
12'd310,  12'd96,  12'd340,  -12'd295,  12'd21,  -12'd204,  -12'd948,  -12'd163,  12'd237,  12'd160,  -12'd55,  12'd510,  12'd43,  -12'd114,  -12'd122,  12'd537,  
12'd145,  -12'd58,  -12'd166,  -12'd186,  -12'd319,  12'd101,  -12'd122,  12'd189,  -12'd231,  -12'd58,  12'd249,  -12'd98,  12'd210,  -12'd61,  -12'd25,  -12'd154,  
-12'd303,  12'd476,  12'd34,  -12'd135,  -12'd74,  12'd297,  -12'd105,  -12'd114,  -12'd238,  12'd172,  -12'd42,  12'd25,  12'd261,  -12'd47,  12'd9,  12'd52,  
12'd69,  -12'd52,  -12'd270,  -12'd87,  12'd49,  -12'd639,  12'd23,  -12'd329,  12'd77,  -12'd171,  -12'd80,  12'd26,  12'd145,  -12'd1,  -12'd214,  12'd416,  
-12'd271,  12'd310,  -12'd229,  12'd51,  12'd361,  12'd168,  -12'd50,  12'd170,  
-12'd198,  12'd409,  -12'd229,  12'd143,  12'd268,  12'd265,  -12'd165,  -12'd109,  -12'd84,  12'd92,  -12'd956,  -12'd118,  12'd288,  12'd59,  12'd338,  12'd467,  
-12'd13,  -12'd80,  -12'd609,  -12'd308,  12'd131,  12'd84,  12'd186,  12'd321,  12'd160,  -12'd405,  -12'd459,  -12'd343,  12'd266,  12'd43,  12'd521,  12'd145,  
12'd86,  12'd292,  12'd376,  12'd311,  -12'd306,  12'd125,  12'd60,  12'd65,  -12'd15,  -12'd209,  12'd357,  -12'd101,  -12'd148,  12'd92,  12'd158,  -12'd559,  
-12'd88,  -12'd300,  -12'd286,  12'd32,  -12'd27,  12'd360,  -12'd301,  12'd387,  12'd219,  12'd339,  -12'd627,  12'd299,  -12'd133,  12'd244,  12'd155,  12'd1,  
12'd149,  -12'd94,  12'd290,  12'd54,  12'd4,  -12'd245,  12'd3,  12'd290,  -12'd132,  -12'd100,  -12'd206,  -12'd171,  12'd74,  12'd312,  -12'd360,  -12'd160,  
12'd170,  -12'd23,  12'd240,  -12'd28,  -12'd622,  -12'd34,  -12'd138,  12'd182,  -12'd306,  -12'd147,  12'd28,  12'd232,  12'd372,  -12'd278,  -12'd365,  -12'd45,  
-12'd19,  -12'd310,  -12'd221,  -12'd73,  -12'd197,  12'd542,  -12'd6,  -12'd355,  -12'd202,  12'd352,  12'd320,  12'd338,  12'd158,  -12'd413,  -12'd180,  12'd58,  
-12'd253,  -12'd153,  12'd105,  -12'd221,  -12'd79,  -12'd23,  12'd171,  12'd302,  
12'd67,  12'd143,  -12'd314,  12'd59,  12'd404,  12'd361,  -12'd83,  -12'd63,  -12'd24,  12'd480,  12'd160,  12'd266,  -12'd5,  12'd97,  -12'd62,  12'd528,  
12'd305,  -12'd152,  -12'd75,  -12'd93,  -12'd31,  -12'd123,  12'd386,  12'd305,  12'd25,  12'd475,  -12'd138,  12'd188,  -12'd161,  12'd237,  12'd230,  -12'd339,  
-12'd222,  -12'd239,  12'd18,  12'd114,  -12'd36,  12'd276,  12'd119,  12'd93,  -12'd438,  12'd193,  -12'd51,  12'd184,  12'd413,  12'd61,  -12'd184,  12'd21,  
-12'd55,  -12'd32,  -12'd179,  12'd399,  12'd385,  12'd520,  12'd315,  12'd380,  -12'd322,  -12'd206,  12'd14,  12'd245,  12'd324,  -12'd60,  12'd183,  12'd43,  
12'd764,  -12'd75,  -12'd89,  -12'd139,  12'd103,  -12'd181,  12'd355,  12'd264,  12'd539,  12'd276,  -12'd385,  12'd122,  -12'd268,  -12'd455,  -12'd120,  12'd19,  
-12'd53,  -12'd292,  -12'd404,  -12'd45,  -12'd31,  12'd224,  12'd42,  12'd54,  -12'd198,  -12'd178,  12'd374,  12'd75,  12'd144,  -12'd463,  -12'd83,  12'd49,  
-12'd38,  -12'd160,  12'd230,  12'd498,  -12'd424,  12'd602,  12'd86,  -12'd113,  12'd116,  12'd240,  12'd321,  12'd155,  -12'd46,  12'd93,  12'd25,  12'd102,  
12'd255,  -12'd50,  12'd62,  -12'd347,  12'd123,  -12'd223,  -12'd162,  -12'd6,  
12'd112,  12'd50,  12'd38,  -12'd32,  12'd146,  12'd182,  -12'd49,  -12'd296,  -12'd208,  12'd108,  -12'd417,  12'd9,  12'd290,  12'd122,  -12'd147,  12'd122,  
12'd197,  12'd402,  -12'd221,  -12'd105,  12'd24,  -12'd183,  12'd332,  -12'd197,  -12'd66,  -12'd550,  12'd4,  -12'd5,  12'd305,  12'd106,  -12'd116,  -12'd36,  
-12'd186,  12'd108,  12'd408,  -12'd131,  -12'd521,  12'd402,  -12'd72,  -12'd350,  12'd131,  -12'd248,  -12'd418,  12'd158,  -12'd124,  12'd18,  12'd347,  12'd283,  
-12'd29,  -12'd633,  12'd316,  -12'd149,  12'd99,  -12'd430,  -12'd20,  -12'd155,  12'd413,  -12'd29,  12'd269,  -12'd21,  -12'd154,  -12'd288,  -12'd234,  -12'd105,  
12'd348,  12'd134,  12'd291,  12'd419,  -12'd196,  -12'd214,  -12'd379,  12'd198,  -12'd289,  12'd328,  12'd181,  12'd284,  12'd281,  12'd351,  -12'd111,  12'd73,  
12'd18,  -12'd143,  -12'd236,  -12'd90,  12'd283,  12'd259,  12'd301,  12'd60,  12'd146,  -12'd21,  12'd329,  12'd229,  -12'd42,  12'd6,  12'd403,  12'd425,  
-12'd210,  12'd75,  12'd175,  12'd240,  -12'd152,  12'd239,  12'd111,  12'd270,  12'd144,  12'd116,  12'd344,  -12'd89,  -12'd124,  -12'd171,  12'd263,  -12'd212,  
12'd53,  -12'd199,  12'd179,  12'd330,  12'd107,  -12'd46,  -12'd315,  12'd27,  
12'd629,  -12'd144,  12'd67,  12'd71,  12'd524,  -12'd273,  -12'd470,  -12'd537,  -12'd5,  -12'd50,  -12'd159,  -12'd292,  12'd160,  12'd168,  12'd96,  12'd222,  
12'd577,  12'd347,  -12'd99,  -12'd42,  -12'd206,  12'd226,  12'd261,  12'd570,  12'd164,  -12'd87,  -12'd204,  -12'd411,  -12'd241,  12'd173,  12'd12,  12'd4,  
12'd442,  -12'd10,  -12'd156,  12'd260,  12'd404,  12'd587,  12'd160,  -12'd285,  12'd79,  12'd229,  -12'd18,  -12'd124,  -12'd96,  -12'd84,  12'd150,  -12'd562,  
12'd4,  12'd144,  -12'd300,  12'd172,  12'd331,  -12'd56,  12'd213,  12'd415,  12'd101,  -12'd28,  -12'd17,  12'd216,  12'd278,  -12'd79,  -12'd242,  -12'd101,  
12'd227,  12'd130,  -12'd192,  12'd26,  -12'd188,  12'd180,  -12'd229,  -12'd356,  12'd184,  -12'd401,  12'd266,  -12'd436,  -12'd78,  12'd34,  -12'd162,  12'd283,  
12'd304,  -12'd2,  -12'd78,  12'd371,  12'd36,  12'd2,  -12'd37,  12'd420,  -12'd83,  12'd43,  12'd310,  -12'd190,  -12'd176,  12'd150,  -12'd207,  12'd80,  
12'd199,  12'd101,  -12'd116,  -12'd388,  -12'd219,  12'd188,  12'd247,  12'd297,  -12'd203,  12'd118,  12'd297,  -12'd416,  12'd298,  12'd377,  -12'd174,  12'd320,  
-12'd344,  -12'd88,  -12'd194,  -12'd15,  -12'd44,  -12'd56,  12'd162,  12'd97,  
12'd49,  -12'd111,  12'd290,  -12'd89,  12'd133,  -12'd100,  12'd174,  -12'd428,  -12'd201,  12'd117,  -12'd371,  -12'd263,  12'd296,  12'd38,  12'd541,  -12'd70,  
12'd290,  12'd199,  -12'd367,  12'd83,  12'd20,  -12'd152,  12'd103,  12'd389,  12'd155,  -12'd63,  12'd71,  -12'd455,  12'd84,  -12'd308,  12'd184,  12'd544,  
12'd257,  -12'd46,  12'd82,  12'd79,  12'd281,  12'd235,  12'd211,  -12'd112,  12'd32,  -12'd234,  -12'd27,  -12'd92,  12'd278,  -12'd341,  -12'd253,  -12'd490,  
-12'd177,  -12'd266,  -12'd222,  12'd539,  -12'd82,  12'd304,  -12'd315,  12'd144,  12'd5,  12'd50,  -12'd293,  12'd369,  -12'd163,  -12'd182,  12'd187,  -12'd202,  
-12'd62,  12'd69,  12'd378,  12'd312,  -12'd86,  -12'd278,  12'd215,  12'd64,  -12'd228,  -12'd152,  -12'd245,  12'd63,  12'd115,  -12'd288,  12'd288,  -12'd133,  
12'd3,  -12'd54,  -12'd216,  12'd208,  12'd5,  -12'd314,  12'd278,  12'd120,  -12'd241,  12'd190,  12'd168,  -12'd90,  12'd316,  12'd45,  12'd97,  -12'd147,  
12'd140,  -12'd90,  -12'd282,  -12'd108,  -12'd188,  12'd554,  12'd170,  12'd7,  -12'd81,  12'd103,  12'd230,  -12'd6,  12'd49,  -12'd299,  -12'd209,  12'd587,  
12'd162,  -12'd134,  -12'd377,  12'd361,  12'd428,  -12'd20,  12'd263,  -12'd87,  
12'd16,  12'd90,  -12'd273,  -12'd106,  -12'd27,  -12'd93,  -12'd30,  -12'd71,  12'd385,  -12'd434,  -12'd3,  -12'd22,  12'd199,  12'd231,  -12'd10,  12'd291,  
12'd26,  -12'd71,  12'd348,  12'd72,  -12'd257,  -12'd51,  -12'd399,  12'd117,  -12'd242,  -12'd310,  -12'd81,  -12'd193,  -12'd173,  12'd146,  -12'd215,  -12'd111,  
12'd207,  12'd173,  12'd77,  -12'd131,  -12'd335,  12'd252,  -12'd243,  -12'd1,  -12'd126,  12'd356,  12'd16,  12'd100,  12'd3,  -12'd98,  -12'd180,  12'd26,  
-12'd21,  12'd7,  12'd127,  -12'd100,  12'd224,  12'd95,  -12'd43,  12'd145,  -12'd127,  12'd21,  -12'd133,  12'd111,  -12'd241,  -12'd181,  -12'd85,  -12'd23,  
-12'd320,  -12'd136,  12'd216,  12'd24,  -12'd288,  -12'd207,  12'd239,  12'd196,  12'd69,  -12'd120,  -12'd146,  12'd234,  12'd1,  -12'd103,  -12'd269,  12'd111,  
12'd387,  12'd175,  -12'd6,  -12'd140,  12'd266,  -12'd210,  12'd79,  12'd231,  12'd49,  12'd193,  12'd27,  -12'd142,  -12'd130,  -12'd21,  12'd189,  -12'd141,  
12'd239,  -12'd327,  12'd149,  12'd54,  -12'd187,  12'd95,  -12'd187,  -12'd155,  -12'd127,  -12'd82,  -12'd106,  -12'd235,  -12'd246,  -12'd109,  12'd74,  12'd67,  
-12'd48,  12'd98,  12'd128,  12'd57,  12'd40,  -12'd115,  -12'd156,  -12'd274,  
-12'd279,  -12'd76,  12'd91,  -12'd84,  -12'd62,  12'd33,  12'd156,  12'd134,  12'd74,  -12'd61,  12'd104,  12'd158,  -12'd221,  -12'd144,  12'd242,  -12'd67,  
-12'd268,  12'd236,  12'd151,  12'd195,  12'd114,  12'd109,  12'd82,  -12'd41,  -12'd162,  12'd136,  12'd45,  -12'd185,  -12'd303,  12'd206,  12'd144,  12'd199,  
-12'd31,  12'd134,  12'd45,  -12'd39,  12'd431,  -12'd99,  -12'd103,  -12'd137,  12'd385,  -12'd281,  12'd136,  12'd125,  12'd271,  12'd203,  12'd185,  12'd274,  
12'd79,  -12'd26,  12'd204,  -12'd166,  12'd53,  12'd463,  -12'd228,  12'd198,  -12'd322,  -12'd52,  -12'd99,  -12'd167,  12'd82,  12'd389,  12'd141,  12'd165,  
-12'd29,  12'd6,  -12'd65,  12'd97,  12'd151,  12'd296,  12'd332,  12'd146,  12'd39,  -12'd315,  12'd116,  -12'd33,  12'd29,  12'd122,  12'd24,  12'd318,  
12'd272,  12'd323,  -12'd70,  12'd395,  12'd197,  -12'd199,  12'd9,  -12'd376,  -12'd88,  -12'd290,  -12'd166,  12'd54,  12'd312,  -12'd243,  12'd29,  -12'd128,  
12'd394,  12'd153,  -12'd205,  -12'd194,  -12'd211,  -12'd392,  12'd90,  -12'd9,  -12'd152,  -12'd182,  -12'd141,  -12'd365,  -12'd69,  12'd110,  -12'd341,  12'd95,  
12'd23,  -12'd36,  12'd128,  12'd125,  -12'd254,  12'd34,  12'd1,  12'd269,  
-12'd284,  12'd180,  12'd18,  -12'd20,  12'd417,  -12'd161,  -12'd36,  -12'd658,  12'd143,  12'd115,  12'd69,  -12'd82,  -12'd106,  -12'd214,  -12'd341,  -12'd333,  
12'd16,  12'd195,  -12'd85,  12'd326,  12'd55,  12'd240,  -12'd387,  12'd234,  12'd106,  12'd80,  12'd490,  12'd83,  12'd152,  12'd79,  12'd151,  -12'd345,  
-12'd116,  -12'd103,  -12'd47,  -12'd202,  -12'd327,  12'd200,  12'd245,  -12'd209,  12'd378,  -12'd52,  -12'd38,  12'd184,  -12'd36,  12'd102,  12'd398,  12'd201,  
12'd14,  12'd30,  -12'd283,  -12'd25,  12'd478,  12'd308,  -12'd496,  12'd99,  -12'd7,  12'd171,  12'd122,  -12'd238,  -12'd5,  12'd334,  12'd23,  -12'd91,  
-12'd94,  -12'd56,  -12'd75,  -12'd174,  12'd115,  12'd139,  12'd47,  -12'd234,  12'd30,  -12'd137,  -12'd64,  12'd61,  12'd388,  -12'd222,  -12'd82,  -12'd22,  
-12'd36,  12'd373,  12'd14,  12'd390,  -12'd243,  -12'd139,  -12'd222,  -12'd54,  12'd126,  12'd224,  12'd278,  -12'd168,  -12'd259,  12'd114,  12'd36,  -12'd225,  
12'd148,  -12'd152,  -12'd369,  12'd137,  -12'd72,  -12'd179,  12'd63,  -12'd744,  -12'd152,  12'd256,  12'd241,  12'd361,  12'd261,  -12'd528,  12'd63,  12'd76,  
12'd108,  -12'd69,  -12'd167,  -12'd195,  12'd51,  -12'd197,  -12'd170,  -12'd292,  
-12'd200,  -12'd18,  12'd329,  -12'd315,  12'd83,  -12'd112,  12'd64,  -12'd206,  12'd100,  12'd304,  12'd251,  -12'd116,  -12'd28,  -12'd8,  12'd163,  12'd275,  
-12'd123,  12'd24,  12'd391,  12'd51,  -12'd95,  12'd284,  12'd59,  -12'd430,  -12'd253,  12'd72,  -12'd188,  -12'd192,  12'd275,  -12'd82,  12'd164,  -12'd305,  
12'd146,  -12'd199,  12'd309,  12'd336,  -12'd401,  -12'd66,  -12'd83,  12'd402,  -12'd340,  -12'd324,  -12'd114,  12'd366,  12'd321,  12'd157,  12'd292,  12'd20,  
-12'd78,  12'd108,  -12'd413,  -12'd370,  -12'd187,  12'd347,  -12'd627,  12'd86,  12'd364,  12'd33,  -12'd76,  12'd155,  -12'd159,  12'd23,  -12'd146,  12'd164,  
12'd84,  12'd331,  -12'd153,  12'd23,  12'd142,  12'd190,  12'd28,  -12'd6,  12'd108,  12'd219,  12'd142,  12'd446,  12'd150,  12'd92,  12'd53,  12'd194,  
12'd75,  -12'd221,  -12'd237,  12'd17,  -12'd187,  -12'd242,  12'd132,  12'd5,  12'd211,  -12'd151,  -12'd86,  -12'd199,  -12'd247,  12'd193,  -12'd100,  -12'd129,  
12'd288,  12'd170,  -12'd162,  12'd440,  12'd124,  -12'd0,  12'd66,  -12'd204,  -12'd70,  12'd231,  -12'd191,  -12'd191,  12'd317,  -12'd466,  12'd233,  -12'd57,  
12'd397,  -12'd36,  12'd148,  12'd18,  12'd67,  -12'd257,  -12'd361,  -12'd13,  
-12'd520,  -12'd33,  -12'd357,  -12'd62,  -12'd153,  12'd167,  12'd157,  -12'd319,  12'd122,  12'd89,  12'd337,  -12'd194,  12'd194,  -12'd194,  12'd132,  -12'd201,  
-12'd230,  -12'd29,  -12'd9,  12'd426,  -12'd176,  -12'd158,  12'd196,  -12'd503,  -12'd141,  12'd24,  12'd11,  12'd513,  12'd181,  -12'd360,  12'd363,  -12'd20,  
12'd65,  -12'd155,  12'd71,  12'd20,  -12'd200,  -12'd1,  -12'd159,  12'd145,  12'd285,  12'd106,  -12'd303,  12'd395,  -12'd389,  12'd2,  12'd443,  -12'd160,  
12'd94,  12'd51,  12'd115,  12'd43,  -12'd29,  12'd54,  -12'd9,  -12'd178,  12'd371,  -12'd367,  12'd347,  -12'd437,  12'd191,  12'd314,  12'd116,  -12'd153,  
12'd33,  12'd132,  -12'd77,  -12'd32,  12'd93,  -12'd218,  12'd320,  12'd98,  -12'd3,  12'd220,  -12'd318,  12'd479,  -12'd269,  12'd435,  -12'd207,  12'd61,  
-12'd153,  12'd14,  12'd242,  12'd185,  -12'd20,  12'd278,  -12'd124,  12'd70,  -12'd22,  12'd213,  -12'd193,  12'd245,  -12'd289,  12'd197,  12'd199,  12'd59,  
-12'd178,  12'd340,  -12'd313,  12'd61,  12'd257,  -12'd133,  -12'd84,  -12'd116,  12'd322,  12'd6,  -12'd57,  12'd89,  -12'd95,  12'd381,  12'd179,  12'd103,  
-12'd3,  -12'd69,  -12'd140,  12'd443,  12'd60,  -12'd382,  12'd334,  -12'd382,  
-12'd153,  -12'd397,  12'd255,  12'd87,  -12'd389,  -12'd101,  -12'd5,  12'd454,  -12'd377,  -12'd278,  -12'd167,  -12'd125,  -12'd317,  -12'd25,  12'd19,  12'd165,  
-12'd85,  -12'd151,  -12'd233,  -12'd35,  -12'd185,  12'd101,  12'd175,  12'd59,  -12'd134,  12'd189,  12'd266,  12'd42,  -12'd271,  -12'd96,  -12'd326,  12'd202,  
12'd70,  12'd359,  -12'd83,  -12'd78,  12'd140,  -12'd46,  -12'd231,  -12'd97,  -12'd52,  12'd74,  12'd324,  -12'd271,  -12'd204,  -12'd234,  12'd154,  -12'd172,  
12'd224,  12'd165,  12'd104,  12'd21,  -12'd532,  -12'd246,  12'd107,  -12'd251,  -12'd270,  12'd389,  12'd9,  -12'd195,  -12'd198,  12'd67,  12'd693,  -12'd116,  
-12'd69,  -12'd493,  -12'd78,  -12'd277,  -12'd106,  -12'd12,  12'd368,  -12'd111,  -12'd132,  12'd80,  -12'd168,  -12'd29,  -12'd128,  12'd284,  12'd6,  12'd215,  
12'd12,  -12'd280,  12'd353,  12'd341,  -12'd166,  12'd224,  -12'd274,  -12'd321,  12'd328,  -12'd107,  -12'd57,  -12'd158,  -12'd153,  12'd32,  12'd207,  12'd108,  
12'd56,  12'd109,  -12'd18,  -12'd33,  12'd363,  12'd505,  12'd122,  -12'd199,  12'd113,  12'd551,  12'd220,  -12'd68,  -12'd120,  12'd760,  -12'd301,  12'd54,  
12'd127,  -12'd429,  12'd271,  -12'd68,  -12'd308,  -12'd320,  -12'd142,  -12'd188,  
12'd121,  -12'd159,  12'd293,  12'd362,  -12'd114,  -12'd115,  -12'd177,  -12'd74,  -12'd41,  12'd414,  12'd112,  12'd57,  -12'd122,  12'd451,  12'd268,  12'd414,  
-12'd101,  12'd185,  12'd95,  -12'd335,  12'd350,  12'd127,  -12'd149,  12'd79,  -12'd353,  12'd60,  12'd93,  12'd135,  -12'd257,  12'd178,  12'd92,  12'd355,  
-12'd110,  12'd40,  12'd91,  -12'd103,  12'd96,  -12'd582,  -12'd288,  12'd35,  -12'd456,  12'd230,  -12'd202,  -12'd202,  12'd447,  12'd217,  12'd148,  -12'd407,  
12'd140,  -12'd34,  -12'd25,  12'd33,  12'd112,  -12'd38,  -12'd245,  -12'd406,  -12'd197,  12'd241,  12'd115,  12'd445,  12'd214,  12'd44,  12'd184,  12'd273,  
12'd175,  12'd188,  12'd153,  -12'd398,  12'd212,  -12'd36,  12'd409,  12'd189,  -12'd124,  -12'd280,  -12'd325,  -12'd102,  12'd396,  -12'd179,  -12'd254,  12'd100,  
12'd294,  -12'd98,  12'd88,  12'd198,  12'd263,  12'd259,  -12'd211,  -12'd150,  -12'd55,  -12'd34,  -12'd106,  -12'd121,  -12'd291,  12'd108,  12'd135,  -12'd34,  
12'd274,  -12'd463,  -12'd146,  -12'd149,  -12'd24,  -12'd311,  12'd220,  -12'd531,  -12'd23,  -12'd413,  -12'd135,  -12'd135,  12'd148,  -12'd37,  -12'd72,  12'd224,  
12'd89,  -12'd259,  -12'd208,  12'd197,  -12'd147,  -12'd404,  12'd160,  12'd47,  
12'd26,  12'd100,  -12'd241,  12'd235,  -12'd151,  12'd341,  12'd38,  -12'd206,  -12'd165,  -12'd377,  -12'd277,  -12'd258,  12'd136,  -12'd90,  -12'd278,  12'd200,  
-12'd78,  12'd91,  -12'd343,  12'd82,  -12'd227,  12'd41,  12'd251,  12'd79,  -12'd57,  12'd181,  -12'd252,  -12'd298,  -12'd86,  -12'd201,  -12'd256,  -12'd2,  
-12'd135,  12'd11,  12'd159,  -12'd233,  -12'd73,  12'd176,  -12'd220,  -12'd218,  12'd169,  -12'd12,  -12'd75,  12'd18,  -12'd152,  12'd64,  -12'd413,  -12'd13,  
12'd208,  -12'd366,  -12'd29,  -12'd270,  -12'd210,  -12'd61,  -12'd113,  -12'd18,  -12'd144,  12'd18,  -12'd302,  12'd33,  -12'd201,  -12'd76,  12'd399,  -12'd141,  
-12'd369,  -12'd328,  -12'd358,  -12'd71,  -12'd169,  -12'd89,  12'd254,  -12'd200,  -12'd188,  12'd77,  -12'd251,  12'd333,  -12'd141,  12'd37,  -12'd290,  12'd80,  
-12'd162,  12'd378,  -12'd55,  -12'd1,  -12'd164,  12'd45,  12'd111,  -12'd93,  12'd119,  -12'd314,  12'd253,  12'd287,  -12'd2,  12'd53,  12'd61,  12'd0,  
-12'd222,  -12'd327,  -12'd24,  -12'd301,  -12'd434,  -12'd17,  -12'd12,  12'd37,  -12'd398,  -12'd169,  -12'd337,  12'd128,  -12'd248,  -12'd73,  12'd49,  -12'd333,  
-12'd393,  12'd252,  -12'd260,  -12'd335,  -12'd29,  -12'd20,  12'd264,  12'd73,  
12'd235,  -12'd101,  -12'd352,  12'd137,  12'd155,  -12'd186,  12'd20,  12'd65,  -12'd142,  12'd140,  12'd301,  -12'd21,  12'd88,  -12'd187,  12'd97,  12'd9,  
-12'd384,  12'd94,  12'd55,  -12'd192,  -12'd68,  -12'd176,  -12'd258,  12'd117,  -12'd56,  -12'd115,  -12'd228,  12'd135,  -12'd100,  -12'd66,  -12'd99,  12'd91,  
12'd3,  -12'd254,  12'd4,  12'd218,  -12'd280,  -12'd74,  12'd46,  -12'd49,  -12'd61,  -12'd131,  -12'd217,  -12'd184,  12'd51,  -12'd91,  -12'd290,  -12'd201,  
-12'd66,  -12'd61,  -12'd204,  -12'd12,  -12'd89,  -12'd147,  12'd177,  12'd58,  12'd27,  -12'd90,  -12'd161,  12'd255,  12'd19,  -12'd215,  12'd212,  -12'd78,  
12'd229,  -12'd469,  12'd32,  -12'd129,  12'd122,  -12'd164,  12'd91,  -12'd178,  -12'd72,  12'd233,  -12'd231,  12'd151,  -12'd18,  -12'd8,  -12'd137,  12'd171,  
-12'd73,  12'd198,  12'd201,  -12'd382,  -12'd308,  -12'd56,  -12'd229,  12'd204,  -12'd5,  -12'd371,  12'd189,  -12'd147,  12'd144,  -12'd29,  12'd297,  -12'd149,  
-12'd216,  -12'd238,  12'd26,  12'd178,  12'd69,  12'd57,  -12'd442,  -12'd263,  -12'd19,  -12'd290,  -12'd128,  -12'd348,  -12'd197,  -12'd84,  12'd58,  -12'd203,  
12'd41,  12'd12,  -12'd329,  -12'd319,  -12'd311,  -12'd197,  -12'd207,  -12'd4,  
-12'd70,  12'd75,  -12'd216,  12'd0,  -12'd259,  12'd294,  12'd71,  12'd40,  -12'd37,  -12'd408,  12'd268,  -12'd63,  -12'd160,  12'd216,  -12'd216,  -12'd41,  
-12'd159,  -12'd201,  -12'd449,  -12'd254,  -12'd201,  -12'd363,  -12'd43,  -12'd59,  -12'd75,  -12'd295,  -12'd246,  -12'd342,  -12'd115,  12'd194,  -12'd88,  -12'd276,  
-12'd98,  -12'd286,  12'd42,  -12'd28,  12'd351,  -12'd281,  -12'd25,  -12'd318,  -12'd346,  -12'd416,  -12'd66,  -12'd148,  -12'd249,  12'd54,  -12'd171,  -12'd62,  
12'd227,  12'd50,  -12'd205,  -12'd322,  12'd52,  12'd97,  -12'd467,  12'd244,  12'd112,  12'd115,  -12'd138,  -12'd111,  -12'd27,  -12'd72,  -12'd31,  -12'd51,  
12'd271,  -12'd280,  -12'd55,  -12'd340,  -12'd169,  -12'd31,  12'd189,  -12'd88,  -12'd109,  -12'd181,  -12'd208,  -12'd196,  -12'd147,  -12'd330,  -12'd203,  -12'd277,  
-12'd254,  -12'd285,  12'd11,  -12'd145,  12'd150,  -12'd196,  12'd40,  12'd45,  -12'd67,  12'd4,  -12'd74,  12'd76,  12'd77,  -12'd82,  12'd26,  -12'd41,  
-12'd502,  -12'd288,  12'd288,  -12'd425,  -12'd221,  -12'd114,  -12'd185,  12'd268,  12'd60,  12'd61,  -12'd36,  -12'd219,  12'd68,  -12'd286,  -12'd263,  -12'd174,  
12'd66,  12'd56,  12'd49,  12'd28,  -12'd51,  12'd99,  12'd71,  -12'd68,  
12'd110,  -12'd141,  -12'd311,  12'd91,  12'd27,  12'd390,  -12'd21,  -12'd66,  -12'd27,  -12'd271,  -12'd0,  12'd28,  -12'd330,  -12'd332,  12'd301,  -12'd156,  
12'd90,  12'd250,  12'd80,  -12'd99,  12'd236,  12'd135,  -12'd234,  -12'd75,  -12'd128,  12'd145,  12'd206,  -12'd148,  -12'd151,  -12'd123,  -12'd142,  12'd115,  
-12'd34,  12'd44,  -12'd210,  -12'd304,  12'd108,  -12'd31,  12'd234,  -12'd87,  -12'd31,  -12'd341,  -12'd132,  -12'd193,  -12'd112,  -12'd40,  -12'd276,  -12'd90,  
12'd186,  12'd20,  -12'd245,  12'd300,  12'd307,  12'd102,  12'd381,  -12'd164,  12'd48,  12'd36,  -12'd179,  -12'd25,  12'd129,  -12'd28,  12'd114,  12'd6,  
-12'd245,  -12'd378,  12'd77,  -12'd365,  -12'd41,  -12'd174,  -12'd70,  -12'd311,  12'd238,  -12'd90,  12'd283,  -12'd213,  12'd227,  12'd238,  -12'd107,  -12'd20,  
12'd123,  12'd296,  12'd15,  -12'd3,  12'd38,  -12'd393,  12'd76,  -12'd169,  12'd98,  12'd146,  -12'd413,  -12'd159,  -12'd45,  -12'd13,  -12'd212,  -12'd108,  
-12'd98,  -12'd171,  -12'd315,  12'd123,  -12'd66,  -12'd145,  -12'd378,  -12'd78,  -12'd332,  12'd179,  -12'd142,  -12'd135,  -12'd158,  -12'd44,  -12'd267,  -12'd197,  
-12'd153,  -12'd177,  12'd211,  -12'd140,  12'd52,  -12'd41,  -12'd68,  -12'd292,  
-12'd188,  -12'd157,  12'd116,  12'd125,  -12'd488,  12'd272,  12'd138,  -12'd16,  12'd186,  -12'd55,  -12'd222,  12'd186,  -12'd9,  12'd288,  12'd372,  -12'd110,  
-12'd685,  -12'd147,  12'd403,  -12'd281,  12'd19,  -12'd324,  12'd205,  12'd8,  12'd151,  -12'd69,  12'd554,  -12'd210,  -12'd631,  12'd137,  -12'd60,  -12'd73,  
-12'd201,  12'd285,  -12'd588,  -12'd183,  12'd82,  12'd501,  12'd437,  -12'd53,  12'd204,  -12'd160,  -12'd168,  -12'd203,  -12'd6,  12'd22,  -12'd52,  12'd183,  
-12'd220,  12'd208,  12'd237,  12'd48,  12'd49,  12'd22,  12'd75,  -12'd89,  12'd248,  12'd303,  12'd22,  -12'd62,  -12'd604,  -12'd0,  12'd444,  -12'd141,  
12'd62,  -12'd373,  12'd246,  12'd140,  12'd347,  -12'd272,  12'd851,  -12'd19,  -12'd429,  12'd68,  -12'd19,  12'd39,  -12'd67,  -12'd195,  -12'd439,  -12'd337,  
12'd143,  12'd167,  12'd58,  -12'd7,  12'd246,  -12'd278,  -12'd204,  -12'd160,  12'd56,  12'd475,  12'd132,  12'd44,  12'd37,  12'd115,  -12'd342,  12'd129,  
12'd247,  -12'd181,  12'd530,  12'd378,  12'd215,  -12'd151,  -12'd346,  12'd334,  12'd206,  12'd477,  -12'd265,  -12'd506,  -12'd183,  12'd23,  -12'd30,  -12'd73,  
12'd227,  12'd156,  12'd392,  12'd357,  -12'd321,  12'd270,  12'd347,  12'd239,  
-12'd334,  -12'd276,  12'd234,  12'd93,  -12'd246,  -12'd416,  -12'd236,  -12'd104,  12'd116,  12'd96,  -12'd113,  12'd213,  12'd15,  -12'd383,  12'd151,  12'd9,  
-12'd87,  -12'd215,  -12'd342,  -12'd304,  -12'd222,  -12'd66,  -12'd116,  -12'd206,  12'd125,  -12'd20,  -12'd150,  12'd33,  -12'd62,  12'd82,  12'd344,  12'd255,  
12'd113,  -12'd150,  -12'd183,  12'd80,  -12'd34,  12'd109,  12'd27,  -12'd75,  -12'd36,  12'd99,  -12'd457,  12'd143,  12'd85,  12'd175,  -12'd53,  -12'd31,  
-12'd150,  12'd193,  -12'd35,  -12'd180,  -12'd154,  12'd177,  -12'd37,  -12'd213,  -12'd286,  12'd25,  -12'd141,  -12'd235,  -12'd59,  -12'd112,  -12'd52,  12'd204,  
-12'd6,  -12'd349,  12'd126,  -12'd40,  -12'd223,  12'd69,  -12'd171,  -12'd25,  12'd156,  -12'd231,  -12'd53,  -12'd99,  12'd57,  12'd12,  -12'd24,  12'd39,  
-12'd37,  -12'd124,  -12'd109,  -12'd255,  -12'd27,  12'd170,  12'd13,  -12'd427,  12'd213,  12'd36,  -12'd40,  12'd140,  -12'd210,  -12'd258,  12'd66,  -12'd80,  
12'd180,  12'd31,  -12'd168,  -12'd97,  -12'd294,  -12'd36,  -12'd174,  12'd72,  -12'd21,  -12'd9,  -12'd182,  -12'd450,  -12'd106,  12'd85,  12'd36,  12'd22,  
-12'd18,  12'd90,  -12'd131,  -12'd64,  -12'd139,  12'd290,  -12'd132,  12'd93,  
12'd587,  12'd43,  12'd113,  -12'd13,  -12'd122,  12'd98,  12'd102,  -12'd339,  12'd293,  -12'd1,  12'd123,  -12'd441,  12'd6,  -12'd295,  -12'd164,  12'd207,  
12'd160,  -12'd140,  12'd77,  12'd104,  12'd173,  12'd305,  12'd43,  12'd462,  12'd162,  12'd234,  12'd7,  12'd208,  -12'd180,  12'd301,  12'd181,  12'd127,  
12'd123,  -12'd254,  12'd211,  12'd279,  12'd10,  12'd328,  12'd397,  -12'd403,  -12'd148,  12'd365,  -12'd364,  -12'd221,  12'd79,  -12'd316,  -12'd394,  -12'd351,  
-12'd78,  -12'd89,  12'd219,  -12'd298,  12'd117,  12'd129,  12'd138,  -12'd61,  -12'd311,  12'd169,  12'd197,  12'd103,  -12'd202,  -12'd30,  -12'd255,  12'd3,  
12'd351,  -12'd522,  12'd344,  12'd114,  -12'd34,  12'd442,  -12'd139,  -12'd237,  -12'd228,  -12'd349,  12'd13,  -12'd433,  -12'd70,  -12'd146,  12'd368,  -12'd95,  
-12'd102,  12'd84,  12'd294,  -12'd7,  -12'd447,  -12'd303,  12'd150,  -12'd227,  -12'd107,  12'd229,  12'd247,  12'd184,  12'd372,  12'd170,  12'd256,  12'd302,  
12'd255,  12'd453,  -12'd348,  -12'd12,  -12'd40,  -12'd270,  12'd190,  12'd721,  12'd36,  -12'd263,  12'd36,  -12'd266,  12'd22,  12'd495,  -12'd276,  12'd84,  
12'd57,  -12'd367,  -12'd246,  -12'd347,  12'd257,  -12'd221,  -12'd164,  -12'd59,  
-12'd366,  -12'd164,  -12'd254,  12'd54,  12'd18,  12'd126,  12'd1,  -12'd14,  -12'd187,  -12'd107,  12'd173,  12'd26,  -12'd203,  12'd236,  -12'd117,  12'd57,  
-12'd215,  -12'd104,  -12'd171,  -12'd3,  12'd275,  -12'd18,  -12'd92,  -12'd64,  12'd64,  12'd60,  12'd244,  12'd245,  12'd160,  -12'd214,  -12'd60,  -12'd568,  
-12'd67,  12'd27,  12'd225,  -12'd168,  12'd156,  12'd94,  -12'd332,  12'd79,  -12'd130,  12'd307,  -12'd40,  12'd16,  -12'd477,  12'd242,  -12'd130,  12'd90,  
12'd213,  -12'd98,  12'd56,  12'd57,  -12'd215,  12'd385,  12'd466,  -12'd53,  12'd116,  -12'd111,  12'd324,  -12'd359,  12'd35,  12'd361,  12'd429,  -12'd250,  
-12'd262,  -12'd15,  12'd67,  -12'd11,  12'd174,  -12'd220,  -12'd103,  -12'd25,  12'd192,  -12'd150,  -12'd308,  12'd69,  -12'd364,  -12'd113,  -12'd278,  12'd131,  
-12'd138,  12'd82,  12'd8,  -12'd265,  12'd88,  12'd217,  12'd86,  -12'd18,  -12'd4,  12'd227,  12'd108,  12'd403,  -12'd413,  -12'd119,  12'd38,  12'd267,  
-12'd117,  12'd142,  -12'd56,  12'd159,  12'd93,  12'd46,  -12'd242,  12'd24,  12'd35,  -12'd13,  -12'd14,  12'd43,  -12'd17,  12'd16,  12'd102,  -12'd470,  
12'd249,  -12'd48,  12'd276,  -12'd114,  12'd350,  12'd217,  12'd112,  12'd97,  
12'd91,  12'd66,  -12'd285,  -12'd43,  12'd590,  -12'd9,  12'd122,  12'd545,  -12'd32,  -12'd104,  12'd185,  12'd297,  -12'd187,  -12'd352,  -12'd118,  -12'd243,  
12'd524,  12'd256,  -12'd241,  12'd108,  12'd90,  -12'd12,  -12'd41,  12'd45,  12'd20,  12'd353,  -12'd155,  12'd3,  -12'd235,  12'd274,  12'd162,  -12'd318,  
12'd106,  -12'd127,  -12'd157,  12'd57,  -12'd1,  -12'd114,  12'd69,  12'd166,  -12'd128,  -12'd182,  12'd458,  -12'd136,  -12'd76,  12'd317,  -12'd199,  12'd139,  
-12'd57,  12'd326,  12'd105,  12'd334,  12'd165,  12'd20,  -12'd187,  -12'd85,  -12'd223,  -12'd100,  -12'd159,  12'd220,  -12'd40,  12'd41,  -12'd60,  12'd160,  
12'd191,  12'd279,  -12'd176,  12'd164,  12'd215,  12'd254,  -12'd190,  12'd86,  12'd178,  12'd94,  12'd194,  -12'd112,  -12'd76,  12'd200,  -12'd232,  12'd113,  
-12'd333,  12'd161,  -12'd181,  12'd555,  12'd263,  -12'd262,  -12'd250,  -12'd216,  -12'd114,  12'd280,  -12'd413,  -12'd116,  12'd167,  12'd337,  -12'd35,  -12'd195,  
12'd110,  -12'd166,  -12'd233,  12'd299,  12'd45,  -12'd284,  -12'd213,  12'd267,  12'd230,  -12'd189,  -12'd315,  12'd337,  -12'd69,  -12'd533,  -12'd5,  -12'd212,  
-12'd126,  12'd495,  -12'd256,  12'd263,  -12'd105,  12'd49,  -12'd49,  -12'd169,  
12'd338,  12'd4,  -12'd174,  12'd85,  -12'd48,  12'd179,  -12'd258,  12'd373,  -12'd138,  -12'd68,  -12'd92,  -12'd295,  -12'd172,  -12'd184,  -12'd324,  12'd354,  
12'd90,  -12'd306,  -12'd72,  -12'd122,  12'd328,  12'd123,  -12'd211,  -12'd149,  -12'd233,  12'd157,  -12'd289,  -12'd119,  -12'd380,  -12'd206,  12'd173,  -12'd179,  
-12'd12,  12'd51,  -12'd0,  -12'd0,  12'd137,  12'd128,  -12'd129,  12'd67,  12'd57,  12'd29,  -12'd260,  12'd75,  -12'd110,  12'd173,  -12'd44,  12'd16,  
-12'd213,  -12'd82,  12'd33,  -12'd119,  -12'd267,  -12'd205,  -12'd289,  -12'd183,  -12'd125,  12'd7,  12'd172,  -12'd165,  12'd150,  12'd304,  -12'd125,  -12'd13,  
-12'd133,  12'd244,  12'd85,  12'd204,  -12'd222,  -12'd27,  12'd212,  -12'd73,  12'd16,  12'd187,  -12'd66,  12'd257,  -12'd53,  12'd106,  -12'd208,  12'd175,  
-12'd312,  -12'd48,  -12'd67,  12'd119,  12'd126,  -12'd185,  -12'd289,  12'd119,  -12'd57,  -12'd149,  -12'd151,  -12'd156,  -12'd9,  -12'd259,  12'd234,  -12'd85,  
12'd139,  12'd17,  -12'd101,  -12'd87,  -12'd0,  -12'd92,  12'd219,  12'd340,  -12'd19,  -12'd357,  -12'd161,  12'd104,  12'd190,  12'd107,  -12'd111,  -12'd108,  
12'd49,  12'd285,  12'd284,  12'd23,  12'd81,  12'd195,  -12'd54,  12'd352,  
12'd586,  12'd44,  -12'd11,  12'd277,  12'd332,  12'd10,  -12'd58,  12'd170,  -12'd363,  -12'd141,  -12'd26,  -12'd272,  12'd3,  -12'd53,  12'd165,  12'd120,  
12'd127,  12'd206,  -12'd393,  12'd224,  -12'd332,  12'd18,  12'd130,  12'd439,  -12'd290,  12'd374,  12'd117,  12'd340,  -12'd290,  12'd146,  -12'd23,  -12'd206,  
-12'd43,  -12'd177,  12'd52,  -12'd70,  12'd211,  12'd253,  12'd435,  -12'd12,  12'd341,  -12'd51,  -12'd302,  -12'd408,  -12'd263,  -12'd50,  -12'd342,  12'd122,  
-12'd63,  12'd35,  -12'd292,  -12'd236,  12'd346,  12'd115,  -12'd96,  -12'd249,  12'd403,  12'd439,  -12'd35,  -12'd88,  12'd198,  12'd6,  -12'd425,  12'd1,  
12'd29,  12'd339,  12'd334,  12'd187,  12'd250,  12'd134,  12'd17,  -12'd61,  -12'd121,  12'd481,  -12'd177,  -12'd136,  12'd385,  12'd312,  -12'd48,  12'd81,  
-12'd302,  12'd274,  -12'd76,  12'd26,  -12'd120,  12'd190,  -12'd140,  -12'd7,  -12'd9,  12'd345,  -12'd48,  12'd258,  12'd453,  -12'd88,  12'd157,  -12'd110,  
12'd52,  -12'd35,  -12'd123,  12'd151,  -12'd274,  12'd89,  12'd361,  12'd346,  -12'd387,  -12'd8,  12'd82,  12'd85,  12'd129,  -12'd117,  12'd372,  12'd222,  
-12'd312,  12'd136,  12'd93,  -12'd80,  -12'd119,  12'd46,  12'd40,  12'd457,  
-12'd560,  -12'd189,  12'd283,  12'd18,  -12'd157,  -12'd263,  12'd146,  12'd544,  12'd55,  12'd61,  -12'd179,  12'd559,  -12'd7,  12'd204,  12'd438,  -12'd257,  
-12'd77,  12'd269,  12'd99,  -12'd342,  12'd102,  -12'd418,  12'd4,  -12'd80,  -12'd116,  -12'd247,  12'd431,  -12'd48,  -12'd7,  12'd367,  -12'd89,  -12'd68,  
-12'd288,  -12'd141,  -12'd96,  12'd87,  -12'd102,  -12'd292,  12'd43,  12'd175,  12'd26,  -12'd239,  12'd363,  12'd112,  12'd104,  12'd77,  12'd50,  12'd504,  
-12'd364,  12'd250,  12'd487,  -12'd686,  -12'd201,  -12'd552,  -12'd305,  12'd179,  -12'd192,  -12'd121,  12'd236,  12'd36,  -12'd201,  12'd7,  12'd19,  12'd146,  
-12'd616,  12'd233,  12'd163,  -12'd356,  12'd98,  -12'd633,  -12'd70,  12'd78,  -12'd24,  -12'd293,  -12'd18,  -12'd114,  12'd563,  -12'd63,  -12'd253,  -12'd49,  
12'd26,  12'd330,  -12'd75,  -12'd266,  -12'd54,  12'd178,  12'd45,  12'd99,  -12'd119,  12'd174,  -12'd167,  12'd320,  12'd58,  -12'd32,  12'd53,  12'd90,  
12'd227,  12'd12,  -12'd55,  -12'd118,  -12'd79,  -12'd602,  -12'd42,  -12'd207,  12'd32,  -12'd367,  -12'd398,  -12'd8,  12'd194,  12'd50,  12'd248,  -12'd99,  
12'd201,  12'd177,  -12'd27,  12'd136,  -12'd10,  12'd43,  -12'd353,  12'd467,  
12'd140,  12'd2,  12'd358,  -12'd157,  -12'd208,  12'd41,  12'd290,  -12'd231,  12'd475,  12'd196,  12'd83,  12'd112,  -12'd28,  -12'd385,  -12'd239,  12'd433,  
12'd220,  12'd3,  12'd366,  12'd206,  -12'd107,  12'd256,  12'd57,  12'd260,  12'd213,  12'd198,  -12'd18,  -12'd117,  -12'd304,  -12'd114,  -12'd484,  -12'd479,  
12'd304,  -12'd155,  -12'd56,  -12'd43,  -12'd295,  12'd419,  12'd477,  -12'd292,  12'd223,  -12'd21,  12'd55,  12'd165,  -12'd267,  -12'd24,  12'd29,  -12'd124,  
12'd100,  -12'd386,  12'd16,  -12'd310,  12'd64,  -12'd65,  12'd33,  12'd105,  -12'd464,  12'd25,  12'd42,  -12'd153,  -12'd147,  -12'd121,  -12'd394,  -12'd142,  
12'd608,  -12'd360,  -12'd105,  12'd230,  12'd465,  12'd204,  -12'd317,  12'd318,  -12'd14,  -12'd58,  12'd264,  12'd246,  -12'd373,  -12'd131,  12'd45,  12'd196,  
-12'd255,  12'd1,  -12'd188,  12'd70,  -12'd171,  12'd105,  -12'd175,  12'd457,  12'd142,  12'd165,  -12'd182,  12'd108,  12'd197,  12'd67,  12'd134,  -12'd125,  
-12'd104,  -12'd132,  -12'd189,  -12'd17,  -12'd331,  -12'd51,  12'd74,  12'd339,  -12'd150,  12'd112,  12'd52,  -12'd358,  12'd273,  12'd88,  12'd125,  -12'd107,  
-12'd303,  -12'd133,  -12'd234,  12'd22,  12'd189,  12'd133,  12'd11,  12'd229,  
12'd134,  -12'd13,  -12'd446,  12'd87,  -12'd347,  12'd98,  12'd68,  12'd171,  -12'd352,  -12'd106,  -12'd98,  12'd20,  -12'd136,  12'd127,  12'd114,  12'd446,  
12'd176,  -12'd169,  12'd256,  -12'd210,  -12'd239,  -12'd237,  -12'd118,  -12'd239,  12'd123,  -12'd375,  12'd68,  12'd75,  -12'd9,  12'd149,  -12'd61,  -12'd376,  
-12'd338,  12'd9,  -12'd346,  12'd146,  12'd239,  -12'd183,  -12'd265,  12'd118,  -12'd337,  -12'd454,  12'd9,  -12'd40,  12'd202,  -12'd35,  -12'd47,  12'd253,  
12'd241,  -12'd555,  12'd97,  -12'd222,  -12'd173,  -12'd268,  12'd79,  12'd135,  -12'd266,  12'd101,  -12'd10,  12'd141,  -12'd14,  -12'd415,  -12'd408,  -12'd30,  
12'd273,  -12'd118,  12'd176,  12'd15,  -12'd283,  12'd43,  12'd199,  -12'd78,  12'd8,  12'd433,  -12'd354,  -12'd302,  12'd179,  -12'd118,  -12'd370,  -12'd13,  
-12'd82,  -12'd247,  12'd279,  -12'd267,  -12'd327,  12'd186,  12'd11,  12'd306,  -12'd418,  -12'd58,  -12'd195,  -12'd150,  12'd227,  -12'd62,  -12'd47,  12'd292,  
12'd113,  -12'd335,  12'd327,  -12'd292,  -12'd62,  -12'd618,  -12'd229,  12'd69,  -12'd62,  -12'd199,  -12'd202,  -12'd130,  12'd81,  12'd187,  -12'd269,  12'd391,  
12'd286,  -12'd112,  12'd195,  -12'd172,  12'd123,  12'd2,  12'd299,  12'd457,  
-12'd237,  -12'd95,  -12'd267,  12'd35,  -12'd195,  -12'd270,  12'd79,  12'd11,  12'd160,  -12'd269,  -12'd194,  12'd157,  12'd40,  -12'd40,  12'd225,  -12'd179,  
-12'd73,  -12'd33,  12'd26,  12'd151,  12'd273,  12'd101,  -12'd12,  12'd18,  -12'd53,  -12'd160,  -12'd17,  -12'd298,  12'd119,  -12'd380,  -12'd177,  -12'd135,  
12'd279,  -12'd433,  -12'd444,  12'd225,  -12'd154,  -12'd402,  -12'd25,  -12'd311,  -12'd67,  12'd226,  -12'd167,  -12'd263,  -12'd226,  12'd10,  -12'd266,  12'd6,  
12'd162,  12'd155,  -12'd183,  -12'd78,  -12'd98,  12'd67,  12'd36,  -12'd125,  12'd202,  12'd66,  12'd55,  -12'd158,  -12'd293,  12'd15,  -12'd62,  12'd287,  
12'd71,  12'd3,  -12'd150,  -12'd46,  -12'd44,  -12'd1,  -12'd29,  12'd58,  12'd11,  -12'd120,  -12'd233,  12'd145,  -12'd168,  -12'd230,  -12'd187,  12'd217,  
12'd246,  -12'd226,  -12'd211,  12'd395,  -12'd255,  12'd143,  -12'd233,  -12'd202,  12'd209,  -12'd306,  12'd83,  -12'd412,  -12'd162,  -12'd2,  -12'd360,  12'd18,  
12'd189,  -12'd243,  -12'd123,  12'd16,  -12'd129,  12'd216,  12'd139,  12'd106,  12'd196,  -12'd73,  12'd171,  12'd59,  12'd212,  -12'd391,  -12'd33,  12'd53,  
-12'd144,  -12'd182,  -12'd97,  -12'd77,  -12'd252,  -12'd91,  12'd226,  -12'd5,  
12'd50,  -12'd194,  -12'd292,  12'd2,  -12'd58,  12'd83,  -12'd89,  -12'd299,  12'd260,  -12'd214,  12'd247,  -12'd204,  12'd163,  -12'd349,  -12'd87,  12'd63,  
-12'd88,  12'd154,  -12'd25,  12'd54,  12'd132,  12'd193,  12'd237,  12'd81,  12'd371,  12'd138,  12'd89,  -12'd94,  -12'd390,  -12'd89,  12'd237,  12'd175,  
12'd445,  12'd220,  12'd56,  -12'd68,  -12'd15,  12'd55,  12'd236,  -12'd203,  12'd232,  12'd298,  -12'd137,  12'd375,  -12'd75,  -12'd293,  -12'd376,  -12'd482,  
-12'd45,  -12'd187,  -12'd111,  12'd454,  12'd129,  12'd69,  12'd347,  12'd179,  -12'd270,  12'd362,  12'd108,  12'd19,  12'd178,  12'd252,  12'd33,  12'd17,  
12'd78,  -12'd355,  12'd91,  12'd736,  12'd93,  12'd42,  12'd107,  12'd273,  12'd379,  -12'd280,  12'd62,  12'd66,  -12'd450,  12'd139,  -12'd238,  -12'd257,  
12'd373,  12'd247,  -12'd121,  -12'd7,  12'd305,  12'd18,  12'd389,  -12'd11,  12'd139,  -12'd209,  12'd124,  -12'd88,  12'd220,  -12'd17,  -12'd138,  12'd275,  
12'd246,  12'd305,  -12'd272,  -12'd83,  -12'd213,  12'd102,  -12'd71,  12'd358,  -12'd397,  12'd36,  12'd149,  -12'd651,  12'd23,  12'd416,  12'd21,  12'd133,  
-12'd139,  -12'd138,  -12'd110,  -12'd75,  12'd229,  -12'd66,  12'd279,  12'd162,  
12'd209,  -12'd102,  12'd184,  -12'd110,  -12'd351,  -12'd103,  12'd142,  12'd202,  12'd35,  -12'd30,  -12'd117,  -12'd128,  -12'd77,  -12'd146,  12'd83,  12'd354,  
-12'd251,  -12'd282,  -12'd161,  -12'd239,  12'd21,  12'd142,  -12'd118,  -12'd70,  12'd4,  12'd48,  -12'd359,  -12'd93,  12'd412,  -12'd239,  -12'd34,  12'd401,  
-12'd122,  12'd265,  -12'd16,  12'd92,  -12'd108,  -12'd210,  -12'd376,  12'd35,  12'd18,  12'd137,  12'd453,  12'd89,  12'd0,  -12'd160,  12'd199,  -12'd153,  
12'd267,  12'd403,  12'd178,  -12'd18,  -12'd169,  -12'd361,  12'd529,  -12'd372,  -12'd2,  12'd314,  12'd190,  -12'd376,  -12'd275,  12'd101,  -12'd131,  -12'd1,  
12'd248,  12'd224,  12'd55,  12'd118,  -12'd5,  -12'd557,  -12'd269,  12'd210,  12'd292,  -12'd558,  12'd368,  -12'd471,  -12'd484,  -12'd231,  -12'd39,  12'd48,  
-12'd29,  12'd235,  12'd90,  -12'd157,  12'd222,  12'd319,  -12'd232,  -12'd81,  12'd116,  12'd60,  -12'd209,  12'd26,  12'd165,  12'd233,  -12'd395,  12'd38,  
12'd119,  12'd453,  -12'd172,  -12'd557,  12'd475,  -12'd263,  -12'd440,  -12'd202,  12'd268,  -12'd185,  12'd66,  -12'd85,  12'd129,  12'd53,  12'd245,  -12'd4,  
-12'd188,  12'd239,  12'd309,  12'd223,  12'd262,  12'd369,  12'd138,  -12'd242,  
-12'd447,  12'd127,  -12'd101,  12'd98,  12'd12,  -12'd130,  12'd283,  -12'd408,  -12'd474,  12'd0,  12'd176,  12'd413,  12'd22,  12'd29,  -12'd11,  12'd116,  
-12'd356,  12'd51,  12'd215,  -12'd40,  -12'd123,  -12'd94,  12'd208,  12'd7,  12'd197,  -12'd458,  -12'd9,  12'd63,  12'd277,  -12'd95,  12'd288,  -12'd56,  
12'd80,  -12'd190,  12'd230,  12'd61,  -12'd417,  12'd41,  12'd240,  12'd326,  -12'd81,  -12'd174,  -12'd189,  -12'd347,  12'd100,  12'd86,  12'd227,  -12'd79,  
-12'd66,  -12'd363,  -12'd243,  12'd198,  -12'd173,  12'd49,  12'd217,  12'd118,  12'd163,  12'd23,  12'd280,  12'd137,  -12'd35,  12'd244,  -12'd32,  -12'd196,  
12'd328,  12'd394,  12'd185,  12'd391,  12'd63,  -12'd350,  -12'd17,  12'd49,  12'd16,  -12'd198,  12'd85,  12'd339,  12'd152,  12'd13,  12'd235,  12'd314,  
12'd162,  12'd113,  12'd120,  -12'd309,  -12'd277,  12'd317,  12'd255,  12'd86,  -12'd139,  12'd297,  12'd30,  12'd65,  -12'd414,  -12'd225,  12'd72,  -12'd17,  
12'd31,  -12'd102,  12'd448,  -12'd270,  12'd82,  12'd137,  -12'd139,  -12'd310,  -12'd55,  12'd295,  12'd86,  -12'd194,  -12'd109,  12'd517,  -12'd179,  -12'd224,  
12'd17,  -12'd463,  12'd174,  12'd75,  12'd215,  12'd236,  12'd437,  12'd303,  
12'd86,  12'd53,  12'd179,  12'd57,  -12'd73,  12'd41,  12'd279,  12'd86,  12'd53,  12'd49,  -12'd167,  12'd84,  12'd223,  12'd89,  -12'd188,  -12'd110,  
-12'd33,  -12'd478,  -12'd39,  -12'd197,  -12'd353,  12'd59,  12'd63,  12'd3,  -12'd76,  -12'd300,  12'd41,  -12'd377,  -12'd269,  12'd114,  12'd282,  -12'd58,  
12'd34,  -12'd315,  -12'd254,  -12'd92,  12'd347,  -12'd273,  -12'd310,  -12'd6,  -12'd205,  12'd24,  12'd190,  -12'd205,  12'd248,  12'd63,  -12'd385,  -12'd322,  
12'd5,  -12'd439,  -12'd401,  12'd121,  12'd100,  -12'd157,  -12'd236,  12'd296,  12'd33,  12'd0,  12'd35,  -12'd171,  -12'd210,  12'd11,  -12'd131,  -12'd302,  
-12'd174,  -12'd48,  -12'd123,  12'd244,  -12'd496,  -12'd99,  -12'd49,  -12'd240,  -12'd242,  -12'd10,  -12'd229,  12'd142,  12'd152,  12'd140,  12'd222,  12'd146,  
-12'd198,  12'd205,  -12'd229,  12'd123,  -12'd426,  -12'd123,  -12'd246,  12'd123,  12'd91,  -12'd110,  -12'd191,  12'd74,  -12'd159,  -12'd110,  -12'd131,  -12'd453,  
-12'd29,  -12'd205,  -12'd57,  -12'd199,  -12'd208,  12'd70,  -12'd374,  -12'd253,  12'd174,  -12'd146,  -12'd201,  12'd212,  12'd128,  12'd277,  -12'd96,  12'd82,  
-12'd12,  12'd87,  12'd98,  12'd11,  12'd291,  12'd154,  -12'd200,  12'd40,  
-12'd330,  -12'd240,  -12'd8,  12'd79,  -12'd175,  -12'd135,  -12'd29,  -12'd106,  12'd255,  -12'd204,  12'd295,  12'd26,  -12'd91,  -12'd138,  12'd257,  -12'd156,  
12'd73,  -12'd82,  -12'd258,  -12'd432,  -12'd125,  -12'd380,  -12'd254,  -12'd449,  -12'd210,  -12'd182,  -12'd44,  -12'd167,  -12'd142,  -12'd352,  -12'd44,  -12'd261,  
-12'd38,  -12'd131,  -12'd13,  -12'd76,  -12'd213,  12'd16,  -12'd37,  -12'd86,  12'd190,  12'd166,  -12'd107,  12'd65,  -12'd230,  -12'd155,  -12'd268,  -12'd56,  
-12'd150,  -12'd388,  12'd11,  12'd6,  -12'd247,  -12'd200,  12'd233,  12'd335,  -12'd42,  12'd324,  12'd103,  -12'd388,  -12'd264,  -12'd234,  -12'd308,  -12'd143,  
-12'd197,  -12'd287,  12'd18,  12'd70,  12'd176,  12'd245,  -12'd33,  -12'd223,  -12'd334,  12'd208,  12'd12,  12'd243,  12'd156,  12'd168,  -12'd256,  -12'd475,  
12'd121,  12'd181,  -12'd329,  12'd153,  -12'd52,  12'd35,  -12'd24,  -12'd409,  -12'd216,  12'd138,  12'd100,  -12'd82,  12'd87,  -12'd415,  12'd158,  12'd141,  
12'd324,  -12'd234,  12'd154,  -12'd204,  -12'd36,  -12'd371,  -12'd183,  -12'd129,  -12'd277,  12'd319,  -12'd46,  -12'd345,  -12'd263,  12'd268,  12'd36,  12'd123,  
-12'd139,  -12'd479,  12'd187,  12'd186,  -12'd344,  -12'd302,  -12'd51,  -12'd147,  
-12'd362,  -12'd47,  -12'd370,  -12'd152,  -12'd337,  -12'd61,  -12'd252,  12'd90,  12'd243,  -12'd263,  12'd96,  12'd34,  -12'd249,  -12'd9,  12'd21,  -12'd435,  
-12'd50,  12'd182,  -12'd435,  12'd95,  -12'd236,  12'd195,  12'd77,  -12'd11,  -12'd88,  12'd223,  12'd175,  12'd24,  12'd45,  12'd203,  12'd413,  -12'd199,  
12'd384,  -12'd38,  -12'd162,  -12'd175,  -12'd61,  -12'd111,  -12'd145,  12'd68,  12'd265,  12'd52,  12'd436,  12'd143,  12'd274,  12'd147,  12'd238,  12'd109,  
-12'd51,  12'd84,  12'd403,  12'd282,  -12'd422,  -12'd34,  12'd16,  -12'd342,  12'd117,  12'd52,  -12'd84,  -12'd74,  -12'd315,  12'd250,  12'd152,  12'd66,  
-12'd293,  12'd101,  -12'd191,  -12'd128,  12'd96,  -12'd240,  12'd10,  -12'd187,  12'd172,  -12'd556,  -12'd68,  -12'd122,  -12'd496,  12'd507,  -12'd184,  12'd399,  
-12'd67,  -12'd80,  12'd224,  -12'd125,  12'd224,  12'd326,  -12'd119,  -12'd174,  -12'd70,  -12'd53,  12'd208,  12'd56,  -12'd88,  12'd207,  12'd34,  -12'd134,  
-12'd71,  12'd193,  -12'd231,  -12'd480,  12'd299,  -12'd251,  -12'd407,  12'd42,  12'd26,  12'd17,  12'd41,  -12'd395,  12'd52,  12'd318,  12'd111,  -12'd245,  
-12'd267,  12'd152,  -12'd248,  -12'd101,  -12'd50,  12'd248,  -12'd37,  12'd27,  
-12'd15,  12'd179,  12'd269,  -12'd358,  -12'd145,  12'd80,  -12'd275,  -12'd359,  -12'd271,  12'd425,  -12'd139,  -12'd354,  12'd428,  12'd129,  12'd36,  -12'd196,  
-12'd12,  12'd282,  -12'd122,  12'd342,  12'd62,  12'd214,  -12'd27,  -12'd645,  -12'd39,  12'd281,  12'd198,  -12'd388,  -12'd32,  -12'd235,  12'd22,  -12'd6,  
-12'd115,  12'd89,  12'd59,  12'd123,  -12'd234,  -12'd327,  -12'd320,  -12'd68,  12'd235,  -12'd79,  -12'd344,  -12'd10,  -12'd115,  12'd21,  12'd31,  -12'd10,  
12'd203,  -12'd245,  12'd85,  -12'd375,  12'd465,  12'd58,  -12'd497,  -12'd124,  12'd50,  12'd557,  12'd178,  12'd20,  12'd445,  -12'd117,  -12'd299,  12'd121,  
-12'd285,  -12'd20,  -12'd80,  12'd235,  12'd224,  -12'd285,  -12'd127,  12'd278,  -12'd444,  -12'd263,  12'd502,  12'd319,  12'd131,  -12'd311,  12'd221,  12'd333,  
12'd151,  -12'd241,  -12'd258,  12'd7,  12'd78,  12'd353,  12'd163,  -12'd144,  12'd121,  -12'd88,  -12'd229,  12'd110,  12'd131,  -12'd158,  -12'd375,  12'd317,  
12'd129,  -12'd33,  -12'd229,  -12'd325,  12'd455,  -12'd41,  12'd29,  12'd39,  -12'd232,  12'd414,  12'd244,  -12'd311,  -12'd133,  -12'd75,  -12'd160,  12'd150,  
12'd53,  -12'd231,  -12'd90,  -12'd121,  12'd392,  -12'd120,  12'd283,  12'd446,  
12'd278,  12'd76,  12'd447,  -12'd101,  12'd179,  12'd125,  12'd260,  -12'd438,  12'd39,  -12'd67,  -12'd60,  -12'd246,  12'd298,  -12'd65,  -12'd391,  12'd253,  
12'd91,  12'd262,  -12'd330,  -12'd179,  12'd145,  12'd5,  12'd267,  12'd400,  -12'd66,  12'd119,  -12'd133,  -12'd155,  -12'd116,  12'd155,  12'd86,  -12'd372,  
-12'd74,  -12'd133,  -12'd261,  -12'd307,  12'd396,  12'd161,  12'd219,  12'd139,  12'd107,  12'd113,  -12'd282,  -12'd318,  12'd121,  -12'd5,  12'd186,  12'd113,  
-12'd270,  -12'd359,  -12'd63,  -12'd131,  -12'd58,  12'd119,  12'd88,  12'd157,  -12'd508,  12'd333,  12'd117,  -12'd147,  12'd312,  12'd129,  -12'd41,  12'd224,  
12'd328,  -12'd293,  12'd469,  12'd81,  -12'd30,  -12'd351,  12'd112,  -12'd128,  12'd247,  12'd123,  -12'd188,  -12'd279,  -12'd269,  -12'd16,  12'd88,  -12'd360,  
12'd54,  12'd220,  -12'd389,  -12'd61,  -12'd57,  -12'd24,  -12'd33,  12'd279,  12'd166,  12'd529,  12'd147,  -12'd95,  -12'd120,  12'd168,  -12'd254,  -12'd1,  
-12'd13,  12'd66,  -12'd101,  -12'd43,  -12'd133,  12'd290,  12'd244,  12'd438,  -12'd166,  12'd318,  12'd5,  -12'd140,  -12'd115,  12'd55,  12'd10,  -12'd66,  
-12'd215,  -12'd563,  12'd268,  12'd5,  12'd16,  -12'd34,  12'd18,  -12'd65,  
-12'd175,  12'd43,  12'd490,  -12'd8,  -12'd276,  -12'd48,  -12'd119,  -12'd196,  12'd34,  -12'd282,  12'd182,  -12'd532,  -12'd207,  -12'd24,  -12'd245,  12'd140,  
-12'd85,  12'd450,  12'd302,  12'd53,  -12'd206,  -12'd280,  12'd46,  12'd0,  12'd354,  12'd69,  12'd416,  12'd49,  -12'd239,  12'd314,  -12'd245,  -12'd387,  
12'd402,  12'd30,  12'd288,  12'd266,  -12'd281,  -12'd66,  12'd58,  12'd145,  12'd191,  -12'd247,  -12'd359,  12'd265,  12'd276,  -12'd155,  -12'd2,  -12'd69,  
12'd328,  12'd6,  12'd119,  -12'd196,  -12'd152,  -12'd41,  -12'd248,  -12'd121,  -12'd329,  -12'd82,  12'd66,  12'd225,  12'd157,  12'd52,  -12'd216,  12'd223,  
-12'd31,  -12'd201,  -12'd96,  -12'd249,  12'd325,  12'd553,  -12'd146,  12'd376,  -12'd296,  -12'd23,  12'd5,  -12'd110,  -12'd184,  -12'd177,  12'd73,  -12'd59,  
12'd239,  -12'd91,  -12'd148,  -12'd64,  12'd141,  -12'd86,  12'd208,  -12'd55,  12'd319,  -12'd214,  12'd33,  -12'd194,  12'd404,  12'd121,  12'd106,  12'd23,  
12'd165,  12'd80,  -12'd44,  12'd150,  -12'd144,  12'd65,  12'd37,  12'd466,  12'd113,  -12'd230,  12'd178,  -12'd302,  -12'd143,  12'd224,  12'd261,  12'd473,  
-12'd141,  -12'd107,  12'd363,  12'd327,  -12'd23,  -12'd170,  -12'd123,  12'd108,  
-12'd8,  12'd188,  12'd121,  -12'd143,  -12'd287,  12'd175,  12'd115,  12'd93,  12'd30,  12'd17,  -12'd40,  -12'd78,  -12'd250,  -12'd187,  -12'd50,  -12'd90,  
12'd161,  -12'd132,  12'd77,  -12'd124,  -12'd34,  -12'd296,  12'd25,  -12'd111,  12'd27,  -12'd315,  -12'd411,  12'd7,  12'd99,  12'd55,  -12'd172,  -12'd221,  
-12'd238,  12'd362,  12'd106,  -12'd182,  -12'd39,  -12'd254,  -12'd143,  -12'd136,  12'd161,  -12'd63,  -12'd44,  -12'd30,  12'd181,  -12'd208,  -12'd136,  12'd94,  
12'd73,  -12'd193,  -12'd118,  12'd131,  12'd82,  -12'd87,  -12'd103,  -12'd226,  -12'd82,  12'd160,  12'd67,  -12'd139,  12'd266,  -12'd267,  -12'd61,  -12'd318,  
-12'd222,  -12'd41,  12'd226,  12'd39,  12'd156,  -12'd23,  -12'd15,  -12'd22,  12'd126,  -12'd116,  12'd229,  12'd25,  -12'd62,  -12'd104,  -12'd81,  -12'd99,  
-12'd45,  -12'd68,  -12'd122,  12'd192,  12'd86,  -12'd318,  -12'd85,  -12'd132,  -12'd177,  12'd225,  -12'd335,  -12'd52,  -12'd153,  -12'd216,  12'd239,  -12'd14,  
12'd264,  12'd12,  12'd42,  12'd40,  -12'd225,  -12'd385,  -12'd35,  -12'd73,  -12'd322,  -12'd76,  -12'd79,  -12'd304,  -12'd82,  12'd22,  -12'd10,  12'd288,  
-12'd190,  -12'd48,  12'd42,  -12'd77,  -12'd225,  12'd103,  12'd15,  -12'd289,  
12'd8,  -12'd34,  -12'd75,  12'd239,  12'd55,  -12'd132,  -12'd321,  12'd115,  -12'd341,  -12'd162,  12'd1,  -12'd302,  -12'd90,  -12'd145,  12'd30,  12'd3,  
-12'd57,  -12'd212,  -12'd190,  12'd68,  -12'd70,  -12'd19,  -12'd31,  -12'd330,  -12'd19,  12'd129,  12'd201,  -12'd203,  12'd109,  -12'd209,  -12'd9,  12'd9,  
12'd90,  -12'd424,  -12'd31,  -12'd300,  -12'd297,  12'd32,  12'd163,  -12'd68,  -12'd264,  -12'd249,  12'd113,  -12'd9,  -12'd8,  -12'd145,  -12'd128,  -12'd18,  
12'd198,  12'd255,  -12'd148,  12'd309,  -12'd129,  -12'd383,  -12'd76,  -12'd22,  -12'd343,  12'd59,  12'd84,  -12'd404,  -12'd42,  -12'd158,  12'd350,  -12'd131,  
-12'd367,  -12'd285,  12'd151,  -12'd64,  -12'd128,  -12'd207,  12'd241,  -12'd174,  -12'd273,  -12'd72,  -12'd150,  -12'd34,  -12'd89,  -12'd407,  12'd86,  -12'd7,  
-12'd94,  -12'd46,  12'd140,  -12'd256,  -12'd204,  12'd151,  -12'd168,  -12'd341,  -12'd338,  -12'd340,  -12'd108,  -12'd148,  -12'd158,  12'd184,  12'd383,  -12'd9,  
12'd139,  -12'd169,  -12'd345,  -12'd25,  12'd274,  12'd203,  12'd267,  12'd107,  -12'd42,  12'd35,  -12'd46,  -12'd135,  12'd85,  12'd26,  -12'd426,  -12'd208,  
-12'd411,  -12'd382,  12'd99,  -12'd352,  -12'd168,  12'd77,  12'd74,  -12'd138,  
12'd9,  -12'd349,  -12'd295,  12'd192,  -12'd55,  12'd73,  -12'd62,  -12'd801,  -12'd372,  -12'd179,  -12'd116,  12'd293,  -12'd40,  12'd101,  12'd213,  -12'd100,  
-12'd104,  -12'd64,  -12'd159,  -12'd73,  12'd70,  12'd108,  12'd241,  -12'd304,  -12'd148,  12'd465,  12'd383,  12'd309,  -12'd93,  12'd217,  12'd213,  12'd281,  
12'd129,  12'd441,  12'd267,  12'd156,  12'd168,  -12'd118,  12'd229,  -12'd206,  12'd229,  12'd362,  12'd26,  -12'd319,  -12'd435,  12'd191,  -12'd145,  -12'd432,  
12'd205,  -12'd208,  12'd74,  -12'd320,  12'd317,  12'd281,  12'd32,  -12'd10,  -12'd198,  12'd54,  12'd169,  12'd118,  12'd198,  -12'd56,  12'd203,  -12'd325,  
12'd85,  12'd208,  -12'd140,  -12'd540,  -12'd56,  -12'd46,  12'd482,  -12'd162,  -12'd49,  -12'd216,  -12'd84,  -12'd275,  12'd103,  -12'd15,  -12'd238,  -12'd138,  
12'd290,  12'd86,  -12'd271,  -12'd308,  12'd265,  -12'd184,  -12'd354,  -12'd265,  -12'd147,  12'd530,  12'd60,  12'd310,  12'd103,  -12'd178,  -12'd268,  12'd102,  
-12'd179,  -12'd147,  -12'd65,  -12'd54,  -12'd46,  -12'd446,  -12'd128,  -12'd286,  12'd131,  -12'd103,  12'd386,  -12'd133,  12'd68,  12'd747,  -12'd24,  12'd264,  
-12'd176,  12'd135,  12'd505,  -12'd38,  -12'd29,  12'd137,  12'd89,  12'd9,  
12'd247,  -12'd53,  12'd213,  12'd194,  -12'd60,  -12'd345,  -12'd62,  12'd29,  -12'd123,  12'd340,  12'd559,  12'd225,  -12'd374,  -12'd303,  -12'd326,  12'd51,  
-12'd173,  -12'd136,  12'd251,  12'd3,  -12'd76,  -12'd237,  12'd281,  12'd232,  -12'd260,  12'd65,  12'd138,  12'd327,  -12'd406,  -12'd82,  12'd97,  12'd30,  
12'd30,  -12'd13,  12'd104,  12'd126,  12'd29,  12'd225,  12'd55,  12'd51,  -12'd53,  12'd98,  12'd179,  -12'd134,  -12'd395,  12'd13,  -12'd706,  -12'd170,  
-12'd175,  12'd243,  -12'd3,  12'd423,  -12'd527,  12'd111,  12'd376,  12'd251,  12'd321,  -12'd466,  -12'd270,  -12'd380,  12'd302,  -12'd246,  12'd205,  12'd130,  
12'd116,  -12'd85,  12'd85,  12'd361,  12'd77,  12'd170,  12'd293,  12'd142,  12'd45,  -12'd331,  -12'd278,  -12'd106,  -12'd403,  -12'd588,  -12'd73,  -12'd86,  
12'd190,  12'd13,  -12'd152,  -12'd357,  12'd477,  12'd49,  12'd19,  -12'd85,  12'd166,  12'd21,  12'd411,  12'd166,  12'd27,  -12'd4,  -12'd314,  12'd30,  
12'd98,  -12'd89,  12'd467,  12'd605,  -12'd165,  12'd665,  -12'd60,  -12'd127,  12'd122,  -12'd110,  12'd125,  12'd118,  12'd78,  -12'd500,  12'd199,  12'd154,  
12'd42,  -12'd214,  12'd143,  -12'd243,  -12'd81,  -12'd177,  12'd221,  -12'd129,  
-12'd36,  12'd146,  12'd87,  -12'd126,  12'd184,  -12'd176,  -12'd0,  12'd404,  12'd604,  -12'd301,  12'd167,  -12'd260,  -12'd321,  -12'd410,  -12'd172,  -12'd50,  
12'd187,  -12'd79,  -12'd145,  12'd379,  -12'd33,  12'd111,  -12'd99,  -12'd85,  12'd7,  12'd112,  -12'd187,  -12'd218,  -12'd299,  12'd79,  12'd464,  12'd154,  
12'd66,  -12'd281,  -12'd155,  12'd152,  12'd522,  12'd130,  12'd16,  12'd345,  12'd44,  12'd13,  12'd218,  -12'd310,  12'd134,  12'd140,  -12'd5,  12'd59,  
-12'd102,  12'd143,  12'd3,  -12'd121,  12'd198,  -12'd7,  12'd6,  12'd112,  12'd63,  -12'd299,  -12'd391,  -12'd148,  12'd235,  12'd89,  12'd186,  12'd95,  
-12'd235,  12'd144,  -12'd70,  -12'd5,  -12'd116,  12'd223,  -12'd67,  12'd53,  12'd416,  -12'd268,  -12'd299,  -12'd452,  -12'd27,  12'd322,  12'd196,  12'd382,  
12'd273,  12'd193,  -12'd173,  12'd502,  -12'd39,  12'd96,  -12'd23,  12'd294,  12'd329,  12'd73,  -12'd231,  12'd245,  12'd378,  -12'd142,  -12'd67,  -12'd61,  
-12'd79,  12'd153,  -12'd756,  -12'd323,  12'd132,  -12'd247,  -12'd494,  12'd553,  12'd237,  -12'd247,  -12'd187,  -12'd232,  -12'd29,  -12'd330,  12'd66,  -12'd82,  
-12'd186,  12'd568,  12'd241,  -12'd138,  -12'd123,  -12'd267,  12'd15,  12'd96,  
12'd32,  -12'd148,  -12'd478,  12'd141,  12'd280,  12'd108,  -12'd62,  -12'd250,  -12'd51,  12'd430,  -12'd513,  12'd143,  12'd158,  12'd139,  12'd318,  -12'd249,  
12'd370,  12'd134,  12'd255,  12'd379,  12'd364,  12'd283,  12'd241,  12'd65,  12'd51,  -12'd394,  -12'd117,  12'd2,  12'd222,  -12'd149,  12'd381,  -12'd312,  
-12'd329,  -12'd297,  12'd243,  12'd61,  -12'd303,  -12'd100,  12'd64,  12'd150,  12'd433,  -12'd318,  -12'd117,  12'd99,  12'd105,  12'd332,  12'd321,  12'd417,  
12'd61,  -12'd315,  12'd249,  -12'd266,  12'd39,  -12'd14,  -12'd385,  12'd80,  12'd54,  12'd76,  -12'd0,  12'd152,  -12'd116,  12'd50,  -12'd410,  12'd179,  
-12'd261,  12'd108,  12'd86,  12'd117,  12'd226,  -12'd295,  -12'd96,  -12'd293,  -12'd267,  12'd233,  -12'd279,  12'd423,  12'd529,  12'd317,  -12'd107,  -12'd26,  
-12'd139,  12'd45,  -12'd267,  -12'd234,  -12'd218,  12'd195,  12'd151,  12'd203,  12'd108,  -12'd129,  -12'd122,  12'd162,  12'd375,  12'd389,  12'd25,  -12'd84,  
12'd317,  -12'd398,  12'd214,  -12'd350,  -12'd3,  12'd94,  -12'd304,  -12'd357,  12'd76,  12'd28,  -12'd380,  12'd307,  -12'd107,  -12'd554,  12'd161,  12'd275,  
-12'd161,  12'd111,  -12'd167,  12'd310,  12'd290,  12'd26,  -12'd201,  -12'd215,  
-12'd364,  -12'd104,  -12'd194,  -12'd13,  -12'd66,  -12'd170,  12'd348,  -12'd460,  12'd563,  12'd172,  12'd234,  -12'd186,  -12'd79,  12'd270,  -12'd115,  12'd235,  
12'd171,  -12'd192,  12'd340,  12'd221,  12'd18,  12'd323,  12'd387,  -12'd392,  -12'd334,  -12'd126,  -12'd214,  -12'd253,  12'd419,  -12'd172,  -12'd287,  12'd490,  
12'd325,  -12'd12,  12'd90,  12'd187,  -12'd281,  12'd150,  12'd96,  -12'd108,  -12'd148,  12'd287,  12'd401,  12'd162,  -12'd96,  12'd90,  -12'd204,  -12'd31,  
-12'd207,  12'd74,  -12'd124,  12'd143,  -12'd43,  -12'd147,  12'd83,  12'd29,  12'd184,  -12'd104,  12'd43,  12'd538,  -12'd89,  -12'd192,  12'd58,  12'd60,  
12'd3,  -12'd196,  -12'd35,  12'd294,  12'd201,  12'd504,  -12'd160,  12'd261,  12'd272,  -12'd275,  12'd275,  -12'd361,  12'd153,  12'd75,  12'd314,  12'd340,  
-12'd258,  -12'd61,  12'd215,  12'd584,  -12'd8,  -12'd127,  12'd246,  -12'd355,  12'd335,  -12'd523,  -12'd339,  -12'd58,  12'd89,  12'd153,  12'd164,  -12'd141,  
12'd236,  12'd223,  -12'd418,  -12'd47,  -12'd174,  12'd75,  12'd20,  -12'd78,  12'd106,  12'd484,  -12'd38,  -12'd420,  12'd56,  12'd75,  -12'd264,  -12'd33,  
12'd150,  12'd327,  -12'd24,  -12'd146,  12'd38,  -12'd382,  12'd36,  -12'd322,  
12'd215,  12'd107,  12'd385,  12'd104,  -12'd132,  12'd76,  12'd257,  12'd590,  -12'd43,  12'd322,  -12'd300,  -12'd110,  -12'd128,  -12'd29,  -12'd247,  -12'd465,  
-12'd378,  12'd217,  12'd116,  -12'd135,  -12'd173,  -12'd204,  -12'd178,  12'd228,  -12'd125,  -12'd94,  12'd299,  12'd31,  -12'd239,  12'd204,  -12'd95,  -12'd58,  
-12'd142,  -12'd47,  -12'd142,  12'd297,  12'd88,  12'd10,  12'd228,  12'd39,  12'd325,  -12'd74,  12'd81,  -12'd44,  12'd120,  -12'd111,  -12'd79,  12'd238,  
12'd228,  12'd388,  12'd15,  -12'd561,  -12'd394,  -12'd192,  12'd123,  -12'd21,  12'd194,  -12'd79,  12'd401,  12'd54,  12'd111,  12'd143,  12'd246,  12'd209,  
-12'd297,  12'd110,  -12'd370,  -12'd380,  -12'd228,  -12'd229,  -12'd397,  12'd111,  -12'd374,  12'd75,  12'd205,  12'd8,  12'd451,  -12'd108,  12'd64,  12'd122,  
12'd236,  -12'd128,  12'd138,  12'd16,  12'd143,  12'd238,  12'd192,  12'd304,  12'd176,  -12'd103,  12'd326,  -12'd353,  -12'd39,  12'd337,  12'd126,  -12'd94,  
-12'd86,  -12'd45,  12'd215,  -12'd64,  12'd322,  12'd62,  12'd343,  12'd237,  12'd31,  -12'd177,  -12'd168,  -12'd385,  -12'd83,  -12'd523,  -12'd140,  -12'd146,  
12'd136,  -12'd42,  -12'd205,  12'd97,  12'd79,  -12'd251,  12'd80,  12'd249,  
-12'd133,  12'd168,  12'd209,  -12'd47,  -12'd27,  -12'd117,  -12'd53,  12'd168,  -12'd29,  12'd415,  12'd207,  -12'd330,  12'd43,  -12'd227,  12'd113,  -12'd668,  
-12'd66,  12'd262,  12'd32,  -12'd185,  12'd25,  -12'd20,  12'd135,  12'd192,  -12'd163,  -12'd92,  -12'd247,  -12'd663,  -12'd18,  -12'd197,  12'd244,  12'd187,  
-12'd140,  12'd238,  -12'd139,  12'd193,  12'd37,  -12'd732,  -12'd220,  -12'd174,  -12'd45,  -12'd321,  12'd245,  -12'd38,  12'd261,  12'd404,  -12'd14,  12'd161,  
12'd133,  12'd220,  12'd161,  -12'd152,  -12'd348,  -12'd346,  -12'd365,  12'd76,  -12'd103,  12'd310,  12'd211,  -12'd59,  -12'd440,  -12'd132,  -12'd268,  12'd23,  
12'd165,  12'd206,  -12'd16,  12'd165,  -12'd153,  12'd41,  12'd344,  -12'd97,  -12'd312,  -12'd405,  12'd96,  12'd192,  12'd225,  12'd347,  12'd20,  -12'd129,  
12'd53,  12'd66,  12'd308,  12'd290,  12'd105,  -12'd3,  -12'd463,  -12'd258,  12'd64,  -12'd309,  12'd170,  -12'd63,  -12'd30,  12'd318,  12'd15,  -12'd328,  
12'd422,  -12'd100,  12'd346,  -12'd153,  12'd13,  12'd11,  -12'd85,  12'd313,  12'd79,  12'd3,  -12'd214,  -12'd665,  -12'd35,  -12'd158,  -12'd564,  12'd304,  
-12'd178,  12'd307,  -12'd481,  -12'd109,  -12'd272,  -12'd151,  12'd215,  12'd197,  
-12'd18,  12'd254,  12'd100,  12'd14,  12'd227,  -12'd78,  -12'd112,  12'd585,  12'd323,  -12'd132,  12'd9,  -12'd52,  12'd0,  12'd34,  12'd409,  12'd98,  
12'd19,  -12'd131,  -12'd167,  12'd347,  12'd351,  12'd99,  12'd266,  12'd41,  12'd161,  -12'd43,  -12'd42,  -12'd35,  12'd276,  12'd402,  12'd256,  12'd299,  
-12'd192,  -12'd73,  -12'd84,  12'd222,  -12'd345,  12'd207,  12'd14,  12'd363,  -12'd296,  -12'd140,  12'd405,  12'd115,  -12'd2,  12'd125,  12'd9,  12'd318,  
-12'd368,  12'd56,  -12'd4,  12'd291,  -12'd197,  12'd13,  -12'd192,  -12'd16,  12'd115,  -12'd554,  -12'd84,  12'd285,  -12'd243,  12'd439,  12'd154,  12'd51,  
-12'd217,  -12'd138,  -12'd27,  12'd148,  12'd34,  -12'd55,  -12'd90,  -12'd133,  12'd165,  -12'd42,  -12'd12,  12'd14,  12'd148,  -12'd1,  -12'd92,  -12'd269,  
-12'd274,  12'd85,  12'd238,  12'd28,  -12'd39,  12'd66,  -12'd67,  -12'd130,  12'd195,  -12'd136,  12'd128,  12'd134,  -12'd6,  12'd3,  12'd112,  -12'd75,  
12'd94,  12'd261,  -12'd655,  12'd119,  -12'd6,  -12'd171,  -12'd357,  -12'd237,  12'd15,  12'd138,  12'd19,  -12'd62,  -12'd119,  -12'd298,  -12'd378,  -12'd4,  
12'd250,  12'd538,  -12'd94,  12'd82,  -12'd215,  12'd56,  12'd137,  -12'd293,  
-12'd202,  12'd146,  -12'd344,  12'd68,  -12'd28,  12'd64,  -12'd238,  -12'd671,  -12'd508,  -12'd318,  -12'd73,  -12'd300,  -12'd437,  -12'd42,  -12'd198,  -12'd25,  
-12'd256,  -12'd222,  -12'd19,  -12'd185,  -12'd246,  -12'd94,  -12'd29,  12'd99,  -12'd32,  -12'd204,  -12'd258,  -12'd26,  -12'd105,  -12'd218,  -12'd137,  -12'd6,  
-12'd59,  12'd296,  12'd243,  -12'd179,  12'd152,  -12'd90,  -12'd199,  12'd232,  -12'd175,  12'd26,  12'd64,  12'd237,  12'd130,  -12'd44,  -12'd139,  -12'd292,  
-12'd97,  -12'd63,  12'd139,  12'd156,  12'd72,  -12'd244,  12'd156,  -12'd177,  -12'd125,  -12'd387,  -12'd183,  -12'd334,  -12'd424,  -12'd134,  12'd18,  -12'd22,  
-12'd147,  12'd85,  12'd143,  12'd286,  12'd1,  -12'd97,  12'd461,  -12'd334,  12'd75,  -12'd207,  12'd249,  -12'd144,  -12'd201,  -12'd392,  -12'd369,  -12'd234,  
12'd3,  -12'd191,  12'd2,  -12'd247,  -12'd249,  -12'd260,  12'd165,  12'd73,  -12'd250,  -12'd110,  12'd121,  12'd111,  12'd91,  -12'd39,  12'd129,  -12'd196,  
-12'd413,  -12'd113,  12'd276,  12'd298,  12'd243,  -12'd21,  -12'd331,  -12'd460,  12'd38,  -12'd308,  -12'd143,  -12'd280,  12'd139,  -12'd130,  -12'd38,  -12'd274,  
-12'd10,  12'd65,  -12'd7,  12'd19,  -12'd92,  12'd30,  -12'd0,  -12'd300,  
-12'd15,  12'd240,  12'd89,  -12'd238,  12'd16,  -12'd179,  12'd109,  -12'd87,  12'd62,  12'd13,  12'd248,  -12'd176,  -12'd215,  -12'd179,  -12'd59,  -12'd5,  
12'd456,  12'd171,  -12'd16,  12'd333,  -12'd144,  12'd198,  -12'd58,  -12'd723,  12'd60,  -12'd166,  12'd176,  12'd269,  -12'd61,  -12'd47,  12'd294,  -12'd220,  
12'd71,  12'd133,  -12'd262,  12'd265,  -12'd248,  12'd246,  -12'd46,  12'd39,  -12'd407,  12'd292,  -12'd37,  12'd207,  -12'd294,  12'd338,  12'd16,  12'd36,  
12'd142,  12'd336,  12'd349,  -12'd82,  -12'd45,  12'd57,  12'd437,  -12'd224,  12'd245,  -12'd311,  -12'd189,  -12'd485,  12'd54,  12'd98,  12'd117,  -12'd326,  
-12'd240,  12'd348,  12'd67,  12'd106,  -12'd55,  -12'd377,  12'd97,  12'd117,  12'd425,  -12'd174,  12'd74,  -12'd235,  -12'd540,  -12'd75,  -12'd422,  -12'd103,  
12'd149,  -12'd10,  12'd136,  -12'd54,  12'd466,  12'd343,  12'd146,  -12'd148,  -12'd265,  -12'd416,  12'd3,  12'd250,  -12'd180,  12'd70,  12'd23,  -12'd173,  
12'd103,  -12'd69,  -12'd146,  12'd9,  12'd366,  12'd144,  -12'd222,  -12'd203,  12'd373,  -12'd165,  12'd35,  12'd149,  -12'd149,  12'd637,  -12'd199,  -12'd186,  
12'd61,  12'd324,  -12'd7,  -12'd341,  -12'd186,  12'd221,  12'd65,  -12'd15,  
-12'd357,  12'd22,  -12'd308,  12'd163,  12'd113,  12'd290,  12'd45,  12'd244,  -12'd415,  12'd371,  -12'd509,  12'd191,  12'd74,  12'd364,  12'd183,  -12'd428,  
12'd371,  12'd332,  -12'd126,  -12'd208,  -12'd189,  12'd61,  12'd158,  12'd199,  -12'd68,  -12'd3,  -12'd92,  12'd146,  12'd557,  12'd238,  12'd668,  12'd69,  
-12'd109,  12'd355,  12'd91,  12'd98,  12'd57,  -12'd287,  -12'd48,  -12'd40,  12'd139,  -12'd223,  -12'd328,  -12'd316,  -12'd53,  12'd72,  -12'd133,  12'd171,  
-12'd321,  -12'd87,  -12'd10,  -12'd81,  12'd96,  -12'd282,  -12'd557,  12'd160,  12'd65,  12'd340,  12'd112,  12'd136,  -12'd112,  12'd171,  -12'd36,  -12'd58,  
-12'd90,  12'd161,  -12'd226,  -12'd181,  -12'd14,  -12'd283,  -12'd59,  12'd171,  -12'd208,  -12'd72,  -12'd42,  12'd189,  -12'd112,  12'd215,  -12'd263,  12'd161,  
12'd190,  12'd151,  12'd177,  12'd203,  -12'd81,  -12'd238,  -12'd50,  12'd205,  12'd163,  -12'd199,  -12'd456,  12'd351,  -12'd293,  -12'd0,  12'd383,  12'd74,  
12'd195,  -12'd174,  12'd17,  -12'd188,  12'd187,  12'd12,  -12'd252,  -12'd428,  -12'd36,  12'd92,  12'd58,  12'd142,  -12'd114,  -12'd211,  12'd78,  -12'd275,  
12'd533,  -12'd134,  -12'd294,  12'd10,  12'd218,  -12'd256,  12'd58,  -12'd225,  
12'd309,  -12'd11,  12'd352,  12'd51,  -12'd186,  12'd332,  -12'd350,  12'd211,  -12'd273,  -12'd326,  12'd49,  12'd77,  -12'd219,  12'd43,  12'd107,  -12'd61,  
12'd211,  -12'd180,  12'd195,  12'd197,  -12'd188,  -12'd155,  12'd47,  -12'd15,  -12'd61,  -12'd22,  12'd373,  12'd307,  -12'd389,  -12'd89,  -12'd5,  12'd3,  
-12'd64,  -12'd153,  12'd18,  12'd233,  12'd283,  -12'd203,  12'd63,  -12'd308,  12'd313,  12'd405,  12'd464,  -12'd136,  -12'd75,  -12'd317,  12'd69,  -12'd257,  
12'd15,  12'd58,  12'd122,  12'd263,  12'd57,  -12'd24,  12'd149,  -12'd356,  -12'd354,  12'd17,  -12'd193,  -12'd393,  12'd51,  -12'd129,  12'd276,  12'd24,  
12'd41,  12'd339,  12'd127,  -12'd17,  12'd191,  12'd394,  12'd144,  12'd32,  12'd264,  -12'd134,  -12'd118,  12'd87,  -12'd61,  -12'd346,  -12'd493,  -12'd314,  
-12'd167,  12'd172,  -12'd71,  -12'd276,  12'd290,  12'd132,  12'd177,  12'd15,  12'd281,  12'd439,  12'd142,  12'd99,  -12'd150,  12'd379,  -12'd68,  12'd448,  
-12'd121,  -12'd367,  12'd148,  -12'd62,  12'd103,  -12'd233,  12'd89,  12'd516,  12'd94,  -12'd6,  -12'd101,  12'd428,  12'd278,  12'd235,  12'd519,  12'd99,  
-12'd96,  -12'd35,  12'd433,  12'd13,  12'd21,  -12'd326,  -12'd422,  12'd179,  
-12'd397,  12'd185,  -12'd18,  -12'd178,  -12'd167,  12'd327,  12'd156,  -12'd111,  12'd80,  -12'd85,  -12'd284,  -12'd127,  -12'd251,  12'd79,  -12'd117,  12'd9,  
-12'd36,  12'd316,  12'd180,  12'd58,  12'd289,  -12'd302,  -12'd150,  12'd225,  -12'd215,  12'd84,  -12'd101,  -12'd314,  -12'd291,  -12'd37,  12'd19,  12'd241,  
-12'd170,  12'd114,  12'd35,  12'd0,  -12'd51,  -12'd294,  -12'd27,  -12'd212,  12'd93,  12'd20,  -12'd53,  -12'd58,  -12'd94,  -12'd55,  12'd124,  -12'd150,  
12'd55,  -12'd219,  12'd370,  -12'd80,  -12'd117,  -12'd388,  12'd122,  12'd157,  -12'd62,  -12'd199,  12'd211,  -12'd438,  -12'd46,  -12'd51,  -12'd184,  12'd41,  
12'd66,  -12'd92,  -12'd37,  -12'd130,  12'd111,  12'd45,  12'd91,  12'd203,  -12'd32,  12'd265,  -12'd8,  -12'd292,  -12'd71,  -12'd22,  -12'd277,  12'd176,  
12'd74,  -12'd134,  -12'd215,  -12'd110,  -12'd92,  -12'd96,  -12'd82,  12'd79,  12'd1,  -12'd87,  -12'd168,  -12'd239,  -12'd164,  -12'd205,  -12'd12,  12'd27,  
12'd104,  -12'd246,  -12'd351,  12'd251,  -12'd171,  -12'd168,  -12'd172,  -12'd402,  -12'd44,  12'd27,  -12'd45,  -12'd138,  -12'd38,  -12'd86,  -12'd172,  12'd332,  
12'd139,  12'd224,  12'd223,  12'd107,  -12'd180,  12'd61,  12'd108,  -12'd197,  
12'd416,  12'd137,  -12'd389,  -12'd174,  12'd33,  -12'd223,  -12'd14,  12'd179,  -12'd111,  -12'd275,  -12'd562,  -12'd227,  12'd258,  -12'd197,  12'd177,  -12'd2,  
12'd410,  -12'd71,  12'd80,  12'd528,  -12'd314,  12'd179,  12'd388,  12'd578,  12'd15,  -12'd143,  12'd79,  -12'd166,  12'd48,  12'd28,  12'd407,  -12'd37,  
12'd17,  -12'd216,  -12'd255,  12'd248,  -12'd219,  12'd358,  12'd471,  -12'd165,  12'd218,  12'd5,  12'd141,  12'd58,  -12'd237,  -12'd321,  -12'd103,  12'd62,  
12'd86,  -12'd16,  -12'd204,  12'd268,  12'd179,  -12'd316,  -12'd52,  12'd27,  12'd42,  12'd236,  -12'd220,  -12'd382,  -12'd223,  -12'd84,  -12'd434,  12'd62,  
12'd357,  -12'd130,  12'd155,  12'd593,  -12'd362,  12'd89,  -12'd61,  12'd153,  12'd96,  -12'd58,  -12'd165,  -12'd193,  12'd21,  -12'd42,  12'd141,  12'd23,  
-12'd46,  12'd297,  -12'd54,  12'd205,  12'd171,  -12'd138,  12'd298,  -12'd80,  12'd374,  12'd282,  -12'd83,  12'd48,  12'd106,  12'd325,  -12'd245,  12'd205,  
12'd206,  -12'd191,  -12'd1,  12'd412,  12'd61,  -12'd14,  12'd168,  12'd465,  -12'd59,  12'd5,  12'd252,  12'd141,  12'd363,  12'd253,  12'd422,  12'd34,  
-12'd33,  12'd264,  12'd127,  12'd252,  12'd344,  12'd326,  12'd167,  12'd24,  
12'd135,  12'd179,  -12'd414,  12'd168,  12'd113,  12'd194,  12'd16,  12'd202,  12'd138,  12'd68,  -12'd379,  -12'd239,  12'd312,  -12'd372,  12'd23,  12'd221,  
12'd263,  -12'd180,  12'd36,  -12'd288,  12'd73,  12'd27,  12'd320,  12'd236,  12'd337,  -12'd223,  -12'd136,  12'd81,  12'd235,  -12'd98,  12'd209,  12'd131,  
12'd126,  12'd223,  12'd261,  -12'd33,  -12'd381,  -12'd184,  -12'd55,  12'd107,  -12'd57,  -12'd133,  12'd93,  -12'd242,  12'd470,  12'd221,  -12'd150,  -12'd92,  
12'd126,  -12'd37,  12'd153,  -12'd71,  -12'd292,  -12'd274,  -12'd145,  -12'd194,  12'd494,  -12'd129,  -12'd289,  12'd96,  -12'd2,  12'd266,  -12'd109,  12'd5,  
-12'd318,  12'd551,  12'd170,  -12'd56,  12'd26,  -12'd291,  12'd153,  -12'd330,  12'd135,  12'd15,  12'd335,  12'd88,  12'd379,  -12'd6,  12'd296,  -12'd88,  
12'd11,  12'd425,  12'd73,  12'd76,  -12'd373,  -12'd144,  12'd158,  -12'd137,  -12'd214,  -12'd172,  -12'd12,  -12'd77,  -12'd73,  -12'd48,  -12'd94,  12'd243,  
-12'd29,  12'd129,  -12'd2,  -12'd166,  12'd241,  12'd128,  12'd167,  -12'd361,  -12'd325,  12'd265,  12'd447,  -12'd524,  12'd201,  12'd146,  -12'd28,  12'd221,  
-12'd107,  -12'd170,  -12'd13,  12'd226,  -12'd99,  -12'd399,  -12'd44,  12'd25,  
12'd100,  -12'd118,  12'd19,  12'd117,  -12'd284,  -12'd142,  -12'd61,  -12'd127,  12'd15,  -12'd57,  -12'd445,  12'd435,  12'd390,  12'd173,  12'd219,  12'd190,  
-12'd17,  12'd267,  -12'd7,  -12'd102,  12'd73,  -12'd158,  12'd264,  12'd212,  -12'd180,  12'd95,  -12'd62,  -12'd187,  12'd187,  12'd170,  -12'd325,  12'd442,  
12'd44,  12'd93,  12'd100,  12'd232,  12'd406,  -12'd331,  -12'd126,  12'd69,  12'd393,  12'd214,  -12'd269,  12'd118,  -12'd463,  -12'd71,  12'd41,  -12'd474,  
12'd106,  -12'd467,  12'd206,  12'd497,  -12'd392,  12'd314,  12'd276,  -12'd145,  12'd29,  12'd42,  -12'd190,  -12'd192,  12'd155,  -12'd136,  -12'd301,  -12'd204,  
-12'd92,  -12'd21,  12'd203,  -12'd43,  -12'd67,  -12'd274,  -12'd133,  12'd283,  12'd111,  12'd125,  12'd267,  12'd76,  12'd259,  -12'd75,  12'd287,  12'd79,  
-12'd136,  -12'd373,  -12'd17,  -12'd422,  -12'd109,  12'd197,  12'd296,  12'd213,  12'd299,  -12'd4,  12'd194,  12'd201,  -12'd336,  12'd372,  12'd40,  -12'd60,  
12'd63,  -12'd79,  12'd248,  -12'd302,  -12'd72,  -12'd21,  -12'd9,  -12'd286,  12'd234,  12'd42,  12'd613,  12'd32,  -12'd47,  12'd437,  -12'd178,  12'd490,  
12'd399,  -12'd263,  12'd213,  12'd271,  12'd116,  -12'd189,  -12'd112,  -12'd70,  
12'd62,  12'd79,  12'd332,  12'd56,  12'd152,  12'd52,  12'd318,  12'd59,  12'd71,  -12'd43,  12'd165,  -12'd23,  12'd79,  12'd34,  -12'd238,  -12'd10,  
12'd83,  12'd135,  12'd308,  12'd165,  12'd243,  12'd76,  -12'd253,  -12'd358,  12'd87,  12'd5,  -12'd212,  12'd40,  12'd110,  12'd2,  -12'd280,  -12'd160,  
12'd94,  12'd358,  -12'd114,  -12'd200,  12'd250,  -12'd45,  -12'd287,  -12'd215,  -12'd123,  -12'd134,  12'd600,  12'd442,  -12'd52,  12'd115,  12'd102,  -12'd227,  
-12'd27,  12'd429,  12'd125,  12'd326,  -12'd285,  12'd218,  -12'd275,  -12'd52,  12'd30,  -12'd1,  -12'd291,  -12'd178,  12'd245,  -12'd109,  12'd515,  -12'd413,  
-12'd386,  12'd167,  12'd181,  -12'd138,  12'd94,  12'd117,  -12'd71,  -12'd16,  12'd395,  -12'd193,  -12'd2,  12'd429,  -12'd18,  12'd210,  -12'd28,  -12'd263,  
12'd5,  -12'd72,  12'd527,  12'd363,  12'd73,  12'd48,  12'd103,  -12'd320,  -12'd3,  12'd98,  12'd83,  -12'd139,  -12'd181,  12'd299,  -12'd113,  -12'd153,  
12'd119,  -12'd237,  12'd372,  12'd259,  12'd355,  12'd340,  -12'd64,  -12'd62,  -12'd220,  12'd264,  -12'd178,  -12'd171,  -12'd14,  -12'd109,  -12'd331,  12'd461,  
12'd103,  -12'd23,  12'd230,  -12'd86,  -12'd96,  -12'd92,  -12'd145,  -12'd44,  
12'd214,  -12'd8,  -12'd410,  12'd140,  -12'd293,  -12'd107,  12'd231,  -12'd4,  12'd237,  12'd380,  12'd156,  12'd132,  -12'd81,  12'd473,  12'd68,  -12'd635,  
-12'd513,  -12'd16,  -12'd388,  12'd379,  12'd67,  12'd24,  12'd161,  -12'd251,  12'd171,  -12'd80,  12'd466,  -12'd51,  12'd48,  12'd577,  12'd124,  12'd191,  
-12'd176,  -12'd323,  -12'd377,  -12'd350,  12'd257,  -12'd108,  -12'd14,  -12'd75,  12'd236,  12'd102,  -12'd413,  -12'd303,  12'd97,  12'd313,  -12'd260,  12'd403,  
12'd33,  -12'd469,  -12'd47,  -12'd154,  -12'd7,  -12'd337,  -12'd39,  -12'd34,  12'd113,  12'd548,  12'd22,  -12'd131,  12'd266,  12'd64,  -12'd224,  -12'd344,  
12'd316,  -12'd125,  12'd215,  12'd241,  -12'd116,  -12'd109,  -12'd487,  12'd53,  -12'd54,  12'd167,  -12'd129,  12'd387,  12'd322,  -12'd67,  12'd102,  -12'd208,  
-12'd139,  -12'd161,  -12'd67,  12'd229,  12'd48,  12'd30,  -12'd472,  12'd178,  -12'd117,  12'd220,  -12'd228,  12'd283,  12'd175,  -12'd88,  -12'd251,  -12'd263,  
-12'd124,  -12'd143,  -12'd36,  -12'd375,  12'd228,  -12'd618,  12'd326,  12'd613,  12'd137,  -12'd39,  -12'd264,  12'd107,  12'd41,  12'd268,  12'd357,  -12'd291,  
-12'd190,  12'd289,  12'd380,  12'd152,  12'd30,  -12'd366,  -12'd240,  -12'd195,  
12'd12,  12'd54,  -12'd191,  12'd56,  12'd186,  -12'd45,  -12'd488,  -12'd209,  12'd149,  -12'd7,  12'd162,  -12'd98,  -12'd125,  -12'd75,  -12'd97,  -12'd304,  
-12'd378,  12'd185,  -12'd110,  12'd19,  -12'd199,  -12'd138,  12'd32,  12'd118,  12'd117,  -12'd198,  12'd21,  -12'd110,  12'd16,  -12'd105,  -12'd17,  -12'd269,  
12'd163,  -12'd362,  12'd228,  12'd6,  -12'd22,  -12'd291,  12'd43,  -12'd471,  12'd51,  -12'd30,  12'd318,  -12'd337,  -12'd442,  12'd174,  -12'd112,  -12'd77,  
-12'd189,  12'd130,  12'd15,  -12'd226,  -12'd11,  -12'd260,  -12'd178,  -12'd95,  -12'd171,  12'd52,  -12'd370,  -12'd328,  -12'd161,  -12'd359,  -12'd54,  -12'd280,  
-12'd21,  -12'd172,  12'd33,  -12'd372,  12'd16,  -12'd147,  -12'd473,  -12'd202,  -12'd51,  -12'd357,  -12'd124,  -12'd121,  12'd187,  12'd163,  -12'd2,  12'd182,  
-12'd343,  -12'd164,  -12'd476,  -12'd3,  -12'd332,  -12'd232,  -12'd497,  -12'd89,  -12'd42,  12'd29,  -12'd3,  -12'd56,  -12'd248,  -12'd326,  -12'd68,  12'd207,  
-12'd274,  -12'd221,  -12'd154,  12'd10,  -12'd416,  12'd37,  12'd278,  -12'd154,  12'd50,  -12'd270,  -12'd6,  -12'd133,  -12'd276,  -12'd270,  -12'd111,  -12'd75,  
-12'd120,  12'd83,  -12'd22,  -12'd52,  12'd88,  12'd69,  -12'd153,  12'd224,  
12'd592,  -12'd64,  12'd355,  -12'd100,  12'd507,  -12'd89,  -12'd119,  12'd164,  -12'd495,  -12'd57,  -12'd83,  12'd128,  -12'd408,  12'd462,  -12'd39,  -12'd308,  
12'd488,  12'd95,  -12'd42,  12'd84,  12'd65,  -12'd128,  -12'd249,  12'd194,  12'd9,  12'd447,  12'd88,  -12'd390,  -12'd257,  12'd278,  -12'd56,  12'd208,  
-12'd60,  12'd55,  12'd40,  -12'd145,  -12'd10,  12'd307,  12'd70,  12'd63,  12'd267,  12'd168,  12'd442,  -12'd117,  12'd40,  12'd50,  12'd13,  -12'd449,  
12'd139,  -12'd58,  12'd393,  12'd432,  -12'd0,  12'd401,  12'd119,  -12'd28,  12'd17,  -12'd78,  -12'd75,  -12'd36,  12'd245,  12'd59,  -12'd288,  -12'd484,  
12'd66,  -12'd95,  -12'd73,  -12'd418,  -12'd131,  12'd59,  12'd164,  12'd194,  12'd285,  12'd102,  12'd282,  -12'd213,  12'd120,  12'd231,  12'd338,  12'd165,  
-12'd222,  12'd220,  12'd9,  -12'd6,  -12'd27,  -12'd216,  -12'd354,  -12'd190,  -12'd357,  -12'd25,  12'd445,  -12'd14,  -12'd101,  12'd75,  12'd188,  -12'd470,  
-12'd252,  -12'd291,  12'd56,  12'd186,  12'd343,  12'd299,  12'd98,  -12'd58,  12'd185,  12'd95,  12'd154,  12'd10,  12'd302,  -12'd509,  12'd13,  12'd199,  
-12'd151,  12'd466,  -12'd214,  12'd262,  12'd10,  -12'd111,  -12'd114,  12'd65,  
-12'd257,  -12'd160,  -12'd2,  -12'd230,  12'd96,  -12'd132,  12'd210,  12'd17,  12'd162,  -12'd151,  -12'd234,  12'd46,  -12'd31,  -12'd40,  -12'd149,  12'd0,  
-12'd211,  12'd151,  12'd229,  -12'd260,  -12'd169,  12'd128,  -12'd94,  12'd276,  -12'd98,  12'd221,  12'd321,  12'd128,  -12'd43,  12'd263,  -12'd214,  -12'd237,  
12'd57,  -12'd97,  12'd98,  -12'd72,  -12'd165,  12'd224,  12'd322,  -12'd71,  -12'd113,  12'd112,  -12'd237,  12'd355,  -12'd26,  -12'd198,  -12'd35,  12'd332,  
12'd114,  12'd36,  -12'd150,  -12'd543,  12'd41,  -12'd61,  -12'd64,  12'd38,  12'd306,  -12'd310,  -12'd370,  -12'd313,  12'd183,  -12'd52,  -12'd570,  12'd50,  
12'd162,  -12'd354,  12'd1,  12'd348,  12'd393,  12'd26,  12'd26,  12'd252,  12'd189,  12'd63,  12'd45,  12'd236,  -12'd467,  -12'd28,  12'd201,  -12'd198,  
12'd305,  12'd11,  -12'd4,  12'd254,  12'd45,  -12'd378,  12'd194,  12'd352,  -12'd135,  12'd178,  12'd450,  12'd165,  -12'd22,  12'd6,  -12'd153,  12'd214,  
-12'd179,  -12'd42,  -12'd90,  12'd90,  -12'd150,  12'd193,  -12'd179,  12'd630,  12'd34,  12'd215,  -12'd69,  -12'd185,  12'd102,  -12'd337,  -12'd30,  12'd174,  
-12'd249,  12'd83,  -12'd301,  -12'd218,  12'd58,  12'd274,  12'd9,  12'd184,  
-12'd14,  12'd15,  -12'd277,  -12'd375,  12'd273,  12'd493,  12'd25,  -12'd234,  -12'd129,  -12'd314,  12'd68,  12'd152,  12'd156,  12'd347,  12'd136,  12'd286,  
12'd202,  12'd30,  -12'd383,  -12'd383,  12'd64,  -12'd69,  -12'd201,  12'd189,  12'd285,  -12'd433,  -12'd12,  -12'd264,  -12'd198,  12'd237,  12'd129,  12'd21,  
-12'd115,  12'd121,  -12'd204,  12'd33,  12'd17,  12'd94,  -12'd285,  12'd93,  -12'd234,  12'd312,  -12'd98,  -12'd34,  -12'd73,  12'd86,  -12'd146,  -12'd321,  
12'd217,  12'd130,  12'd99,  -12'd575,  -12'd2,  -12'd178,  12'd227,  -12'd128,  -12'd23,  -12'd30,  -12'd232,  -12'd241,  -12'd338,  12'd165,  -12'd124,  12'd148,  
12'd294,  -12'd9,  -12'd179,  12'd42,  12'd126,  -12'd642,  12'd259,  12'd118,  12'd337,  -12'd495,  12'd214,  -12'd60,  12'd55,  -12'd85,  12'd57,  -12'd296,  
12'd20,  12'd129,  12'd224,  -12'd340,  12'd158,  12'd224,  12'd86,  -12'd79,  12'd381,  12'd75,  12'd162,  12'd169,  12'd159,  -12'd131,  -12'd173,  12'd73,  
-12'd86,  -12'd8,  12'd355,  12'd329,  12'd197,  12'd51,  -12'd83,  -12'd172,  -12'd38,  12'd243,  12'd360,  -12'd105,  -12'd249,  -12'd106,  12'd31,  -12'd45,  
12'd16,  12'd40,  -12'd122,  -12'd43,  -12'd133,  -12'd220,  12'd68,  12'd283,  
12'd5,  -12'd7,  12'd21,  -12'd69,  12'd182,  -12'd116,  -12'd472,  12'd283,  -12'd616,  -12'd77,  -12'd380,  -12'd195,  12'd133,  12'd231,  12'd179,  12'd21,  
-12'd243,  12'd365,  -12'd437,  -12'd87,  -12'd273,  -12'd243,  12'd90,  12'd496,  -12'd7,  12'd252,  -12'd35,  -12'd438,  12'd228,  12'd343,  -12'd343,  12'd483,  
-12'd385,  -12'd4,  12'd127,  12'd150,  12'd560,  12'd268,  12'd58,  -12'd140,  12'd114,  12'd61,  -12'd86,  -12'd289,  12'd17,  -12'd346,  -12'd223,  -12'd626,  
12'd215,  -12'd181,  -12'd377,  12'd115,  12'd195,  12'd42,  -12'd405,  12'd5,  -12'd183,  -12'd96,  12'd208,  12'd48,  -12'd83,  12'd267,  -12'd196,  12'd13,  
12'd296,  -12'd96,  -12'd132,  12'd66,  -12'd38,  -12'd296,  12'd150,  -12'd55,  12'd103,  -12'd247,  12'd183,  -12'd55,  -12'd527,  12'd141,  12'd46,  -12'd219,  
-12'd195,  12'd158,  -12'd483,  -12'd19,  -12'd176,  12'd12,  -12'd153,  -12'd137,  -12'd13,  -12'd46,  -12'd51,  -12'd171,  -12'd37,  -12'd230,  -12'd192,  12'd192,  
12'd105,  -12'd157,  -12'd106,  -12'd612,  12'd23,  -12'd6,  -12'd27,  12'd7,  -12'd167,  12'd259,  12'd49,  -12'd457,  -12'd167,  12'd432,  12'd105,  12'd404,  
-12'd191,  -12'd265,  12'd212,  12'd53,  12'd108,  12'd80,  12'd448,  12'd97,  
-12'd197,  -12'd316,  -12'd155,  -12'd100,  12'd139,  12'd10,  12'd38,  12'd17,  -12'd37,  12'd345,  -12'd131,  12'd292,  12'd37,  12'd86,  -12'd251,  12'd83,  
-12'd20,  -12'd32,  12'd3,  -12'd25,  -12'd156,  -12'd217,  -12'd237,  12'd201,  -12'd125,  12'd34,  12'd77,  12'd276,  -12'd40,  -12'd172,  -12'd341,  12'd217,  
-12'd456,  -12'd0,  12'd273,  -12'd48,  -12'd354,  -12'd64,  12'd175,  12'd213,  12'd225,  -12'd248,  12'd354,  12'd351,  -12'd119,  -12'd57,  -12'd210,  12'd135,  
12'd11,  12'd13,  12'd114,  12'd7,  12'd114,  -12'd181,  -12'd55,  -12'd138,  -12'd225,  12'd198,  12'd330,  12'd24,  12'd274,  -12'd123,  12'd34,  -12'd349,  
-12'd58,  12'd40,  12'd87,  12'd15,  12'd105,  -12'd110,  -12'd111,  12'd4,  -12'd152,  12'd623,  12'd2,  12'd27,  12'd25,  -12'd9,  -12'd350,  12'd259,  
12'd3,  -12'd142,  -12'd285,  -12'd225,  -12'd136,  -12'd38,  -12'd382,  12'd339,  -12'd36,  12'd200,  12'd420,  12'd291,  12'd159,  12'd198,  -12'd255,  12'd358,  
-12'd291,  -12'd132,  12'd499,  12'd112,  12'd98,  12'd186,  12'd161,  12'd146,  -12'd400,  -12'd20,  -12'd9,  12'd458,  12'd20,  12'd92,  12'd93,  12'd85,  
12'd122,  -12'd264,  -12'd210,  12'd25,  12'd383,  12'd446,  -12'd88,  -12'd7,  
-12'd293,  -12'd151,  -12'd110,  -12'd58,  12'd343,  -12'd165,  12'd290,  12'd244,  12'd562,  -12'd144,  12'd221,  -12'd108,  12'd63,  12'd189,  12'd426,  12'd104,  
12'd24,  -12'd235,  -12'd11,  -12'd152,  -12'd25,  -12'd68,  12'd143,  12'd210,  -12'd57,  12'd542,  12'd38,  12'd263,  12'd0,  12'd47,  -12'd156,  -12'd356,  
12'd456,  -12'd62,  12'd138,  12'd81,  -12'd340,  12'd41,  -12'd114,  12'd47,  -12'd255,  -12'd96,  12'd245,  12'd9,  12'd521,  12'd120,  -12'd299,  12'd219,  
12'd16,  12'd109,  12'd24,  12'd143,  -12'd336,  12'd288,  -12'd549,  -12'd56,  12'd98,  -12'd468,  12'd121,  -12'd37,  -12'd137,  12'd226,  12'd402,  12'd437,  
12'd141,  12'd187,  12'd126,  -12'd153,  12'd282,  12'd79,  12'd225,  12'd22,  12'd218,  12'd154,  12'd20,  12'd78,  12'd179,  -12'd42,  -12'd212,  12'd38,  
-12'd340,  -12'd14,  12'd334,  12'd486,  12'd165,  12'd313,  12'd0,  -12'd271,  -12'd171,  12'd88,  12'd268,  -12'd129,  12'd371,  12'd161,  -12'd125,  -12'd259,  
-12'd149,  -12'd215,  -12'd156,  12'd561,  -12'd244,  12'd286,  12'd156,  -12'd111,  12'd244,  -12'd224,  -12'd88,  12'd244,  -12'd10,  -12'd291,  -12'd178,  -12'd48,  
12'd196,  12'd447,  -12'd481,  12'd62,  -12'd149,  -12'd252,  12'd115,  -12'd255,  
-12'd11,  -12'd60,  -12'd397,  12'd179,  -12'd125,  12'd157,  12'd163,  -12'd1,  -12'd25,  12'd60,  -12'd104,  12'd21,  -12'd52,  12'd20,  12'd202,  -12'd162,  
-12'd354,  -12'd123,  12'd384,  12'd66,  12'd30,  -12'd188,  -12'd81,  -12'd300,  -12'd291,  -12'd11,  12'd319,  12'd195,  -12'd210,  12'd128,  -12'd141,  -12'd186,  
-12'd498,  12'd381,  -12'd166,  12'd38,  -12'd3,  12'd35,  -12'd119,  12'd36,  12'd307,  -12'd259,  -12'd258,  12'd82,  12'd19,  12'd123,  12'd412,  12'd448,  
12'd301,  -12'd250,  12'd452,  -12'd37,  12'd88,  12'd311,  -12'd98,  12'd1,  -12'd52,  12'd334,  12'd295,  12'd82,  12'd196,  -12'd4,  12'd654,  12'd27,  
-12'd226,  -12'd52,  12'd99,  -12'd29,  12'd95,  -12'd82,  12'd177,  -12'd35,  12'd34,  12'd46,  -12'd366,  12'd346,  12'd89,  -12'd400,  -12'd184,  -12'd207,  
12'd82,  -12'd111,  12'd226,  -12'd230,  -12'd359,  12'd282,  -12'd151,  -12'd133,  12'd194,  12'd438,  12'd96,  12'd341,  -12'd258,  12'd27,  12'd126,  12'd354,  
-12'd23,  -12'd253,  12'd556,  -12'd191,  12'd107,  -12'd78,  -12'd35,  12'd405,  -12'd314,  -12'd96,  -12'd121,  12'd154,  12'd145,  12'd119,  12'd218,  -12'd103,  
12'd73,  -12'd119,  12'd426,  -12'd22,  -12'd18,  12'd83,  12'd31,  -12'd38,  
12'd152,  -12'd281,  12'd201,  -12'd114,  12'd111,  12'd35,  -12'd105,  -12'd29,  12'd126,  12'd29,  -12'd299,  -12'd0,  12'd331,  12'd9,  12'd382,  -12'd19,  
12'd93,  12'd132,  -12'd167,  12'd259,  12'd122,  -12'd41,  12'd335,  12'd529,  12'd68,  12'd265,  -12'd312,  12'd0,  12'd54,  -12'd150,  12'd198,  12'd100,  
-12'd88,  12'd145,  12'd178,  -12'd267,  12'd169,  -12'd229,  12'd48,  12'd194,  -12'd117,  12'd99,  12'd97,  -12'd52,  12'd393,  -12'd283,  -12'd60,  -12'd428,  
12'd161,  12'd280,  -12'd144,  -12'd204,  12'd181,  -12'd158,  -12'd394,  12'd235,  12'd65,  12'd116,  -12'd93,  12'd259,  12'd72,  12'd128,  -12'd496,  12'd156,  
12'd362,  -12'd19,  12'd162,  12'd100,  12'd439,  12'd175,  -12'd218,  -12'd73,  -12'd172,  -12'd214,  12'd266,  -12'd47,  12'd330,  -12'd170,  12'd195,  -12'd46,  
12'd116,  12'd462,  -12'd393,  12'd266,  -12'd560,  -12'd301,  12'd309,  12'd486,  -12'd29,  12'd23,  -12'd277,  12'd48,  12'd417,  -12'd91,  12'd91,  12'd81,  
-12'd21,  12'd118,  -12'd409,  -12'd268,  -12'd361,  -12'd146,  -12'd79,  -12'd470,  12'd239,  12'd292,  12'd67,  12'd21,  12'd51,  12'd100,  -12'd296,  12'd148,  
12'd263,  12'd41,  -12'd364,  -12'd74,  -12'd79,  -12'd99,  12'd140,  12'd304,  
-12'd142,  12'd169,  -12'd221,  12'd181,  12'd170,  12'd242,  -12'd104,  -12'd352,  12'd194,  12'd246,  12'd127,  12'd181,  12'd314,  12'd221,  -12'd251,  12'd70,  
-12'd32,  12'd190,  12'd181,  12'd379,  -12'd33,  12'd269,  -12'd195,  -12'd418,  -12'd288,  12'd361,  -12'd382,  12'd150,  -12'd96,  -12'd242,  -12'd55,  -12'd247,  
12'd106,  12'd341,  -12'd261,  12'd34,  12'd394,  12'd224,  -12'd358,  -12'd122,  -12'd245,  12'd361,  -12'd278,  12'd144,  -12'd111,  12'd200,  12'd73,  12'd25,  
12'd146,  -12'd190,  -12'd54,  12'd283,  12'd11,  12'd322,  -12'd8,  -12'd122,  -12'd27,  -12'd222,  -12'd373,  -12'd83,  12'd138,  12'd102,  12'd527,  -12'd105,  
-12'd131,  -12'd288,  12'd57,  -12'd41,  12'd58,  12'd248,  12'd76,  12'd430,  12'd31,  -12'd185,  -12'd342,  -12'd454,  -12'd263,  -12'd201,  12'd132,  12'd496,  
12'd30,  12'd214,  12'd7,  -12'd199,  12'd92,  12'd352,  -12'd432,  12'd314,  12'd24,  -12'd378,  12'd372,  -12'd334,  12'd276,  -12'd166,  12'd168,  -12'd33,  
-12'd271,  -12'd98,  -12'd122,  12'd168,  -12'd122,  12'd395,  12'd244,  12'd373,  -12'd105,  12'd69,  -12'd254,  12'd92,  12'd87,  -12'd477,  12'd194,  12'd334,  
-12'd406,  12'd365,  12'd188,  12'd177,  -12'd13,  -12'd115,  12'd137,  12'd76,  
-12'd24,  12'd35,  -12'd522,  12'd355,  -12'd99,  -12'd327,  12'd342,  -12'd57,  12'd45,  -12'd28,  12'd266,  12'd130,  12'd80,  12'd23,  -12'd99,  12'd256,  
-12'd113,  12'd155,  12'd229,  12'd197,  -12'd99,  12'd189,  -12'd8,  12'd75,  12'd375,  -12'd29,  12'd422,  12'd188,  12'd44,  12'd157,  12'd140,  -12'd105,  
12'd242,  -12'd0,  -12'd246,  12'd293,  -12'd283,  12'd480,  12'd210,  -12'd305,  12'd228,  12'd76,  12'd96,  12'd174,  -12'd119,  12'd79,  12'd165,  12'd428,  
-12'd73,  -12'd123,  12'd174,  -12'd192,  12'd410,  -12'd28,  12'd480,  12'd178,  12'd156,  12'd338,  -12'd334,  -12'd222,  -12'd126,  12'd399,  12'd60,  -12'd247,  
-12'd93,  -12'd125,  -12'd123,  12'd280,  12'd158,  -12'd26,  12'd60,  12'd116,  12'd154,  12'd476,  -12'd131,  -12'd213,  -12'd5,  12'd52,  -12'd152,  12'd196,  
12'd293,  12'd119,  -12'd284,  12'd397,  12'd104,  -12'd296,  12'd45,  12'd465,  12'd362,  -12'd97,  -12'd49,  12'd205,  -12'd176,  -12'd139,  -12'd81,  -12'd105,  
12'd306,  -12'd32,  -12'd199,  -12'd55,  -12'd108,  12'd7,  -12'd248,  12'd510,  -12'd192,  12'd267,  12'd128,  12'd141,  12'd220,  -12'd162,  12'd364,  -12'd91,  
-12'd183,  12'd51,  -12'd46,  12'd176,  12'd341,  -12'd73,  12'd218,  -12'd95,  
-12'd602,  12'd126,  12'd219,  -12'd42,  -12'd557,  12'd260,  12'd50,  -12'd136,  -12'd396,  -12'd389,  12'd287,  -12'd176,  -12'd300,  12'd19,  12'd164,  12'd126,  
-12'd365,  12'd63,  12'd88,  12'd85,  12'd168,  -12'd83,  12'd81,  -12'd322,  -12'd162,  12'd19,  12'd322,  12'd269,  -12'd43,  12'd250,  -12'd36,  -12'd213,  
-12'd231,  12'd34,  -12'd265,  12'd16,  12'd636,  12'd237,  -12'd452,  12'd46,  12'd57,  12'd118,  12'd49,  -12'd20,  -12'd173,  12'd89,  12'd43,  12'd5,  
12'd103,  -12'd266,  12'd375,  -12'd318,  12'd135,  12'd7,  -12'd119,  12'd26,  -12'd627,  12'd221,  12'd407,  -12'd143,  -12'd176,  -12'd121,  12'd448,  12'd158,  
12'd319,  12'd58,  12'd309,  -12'd186,  -12'd30,  -12'd3,  12'd92,  12'd54,  12'd227,  -12'd604,  12'd142,  12'd181,  -12'd7,  -12'd219,  -12'd81,  -12'd46,  
12'd16,  12'd244,  -12'd157,  -12'd325,  12'd352,  12'd346,  12'd304,  12'd154,  12'd201,  12'd11,  12'd229,  -12'd202,  -12'd2,  -12'd45,  12'd49,  12'd403,  
12'd228,  12'd41,  12'd159,  -12'd395,  12'd170,  -12'd386,  12'd300,  12'd98,  12'd68,  -12'd208,  -12'd105,  -12'd252,  -12'd61,  12'd924,  -12'd319,  12'd112,  
-12'd234,  -12'd102,  -12'd51,  12'd24,  12'd55,  -12'd27,  -12'd262,  12'd397,  
-12'd620,  12'd110,  -12'd136,  -12'd17,  12'd30,  12'd110,  12'd355,  12'd13,  12'd559,  12'd15,  12'd458,  12'd80,  12'd374,  12'd93,  -12'd154,  12'd32,  
-12'd275,  -12'd5,  12'd337,  12'd379,  -12'd198,  12'd407,  -12'd262,  -12'd337,  -12'd153,  -12'd93,  12'd50,  12'd305,  -12'd63,  12'd25,  12'd177,  -12'd330,  
-12'd221,  -12'd118,  -12'd101,  12'd315,  -12'd173,  -12'd26,  12'd170,  -12'd34,  -12'd84,  12'd253,  -12'd346,  -12'd7,  -12'd214,  12'd54,  12'd194,  12'd538,  
-12'd142,  12'd89,  12'd348,  -12'd97,  -12'd182,  -12'd240,  -12'd103,  -12'd117,  -12'd168,  12'd85,  12'd47,  -12'd292,  12'd234,  -12'd54,  12'd314,  12'd55,  
-12'd196,  12'd35,  12'd92,  12'd432,  12'd48,  12'd233,  12'd175,  12'd219,  12'd117,  -12'd265,  12'd24,  12'd59,  -12'd364,  12'd174,  -12'd264,  12'd182,  
12'd209,  12'd118,  -12'd28,  12'd43,  12'd182,  12'd99,  12'd299,  12'd89,  -12'd58,  12'd180,  12'd15,  12'd232,  -12'd70,  12'd64,  -12'd2,  -12'd88,  
12'd64,  12'd225,  -12'd47,  12'd40,  -12'd394,  12'd109,  -12'd158,  12'd414,  -12'd191,  12'd327,  -12'd33,  -12'd186,  -12'd287,  12'd542,  -12'd84,  12'd41,  
-12'd60,  -12'd253,  12'd445,  12'd331,  -12'd188,  12'd109,  -12'd161,  -12'd28,  
12'd233,  -12'd88,  12'd249,  12'd148,  12'd131,  -12'd218,  -12'd171,  -12'd153,  -12'd34,  12'd147,  -12'd52,  -12'd423,  12'd351,  12'd180,  12'd328,  12'd0,  
-12'd44,  12'd92,  -12'd25,  -12'd144,  12'd252,  -12'd10,  -12'd256,  12'd133,  12'd113,  12'd22,  -12'd98,  -12'd239,  12'd266,  12'd223,  12'd316,  12'd406,  
12'd35,  12'd56,  -12'd252,  -12'd59,  12'd315,  12'd110,  12'd452,  -12'd462,  -12'd180,  12'd324,  -12'd104,  -12'd98,  -12'd138,  12'd30,  -12'd370,  -12'd261,  
-12'd74,  12'd206,  12'd46,  12'd9,  12'd402,  12'd251,  -12'd385,  12'd189,  12'd101,  -12'd329,  12'd83,  12'd130,  12'd152,  12'd40,  -12'd211,  -12'd249,  
12'd369,  12'd39,  12'd64,  -12'd85,  -12'd153,  12'd293,  12'd234,  -12'd62,  12'd26,  -12'd200,  12'd133,  -12'd259,  12'd38,  12'd259,  -12'd186,  -12'd6,  
12'd80,  -12'd79,  -12'd243,  12'd571,  12'd290,  -12'd8,  12'd82,  12'd86,  -12'd410,  -12'd100,  -12'd6,  -12'd441,  12'd126,  12'd200,  -12'd190,  -12'd324,  
-12'd101,  12'd125,  -12'd285,  -12'd21,  -12'd285,  12'd203,  -12'd64,  12'd155,  -12'd333,  12'd309,  -12'd31,  12'd359,  -12'd179,  -12'd75,  12'd342,  12'd141,  
-12'd34,  -12'd54,  12'd93,  -12'd9,  -12'd7,  12'd67,  -12'd59,  -12'd10,  
-12'd473,  -12'd342,  12'd464,  -12'd178,  -12'd212,  -12'd202,  -12'd35,  12'd407,  12'd10,  12'd213,  12'd691,  12'd4,  -12'd143,  12'd234,  -12'd328,  12'd302,  
-12'd346,  12'd144,  12'd295,  -12'd276,  -12'd121,  -12'd49,  -12'd2,  12'd61,  12'd282,  12'd177,  12'd147,  12'd163,  -12'd168,  -12'd86,  -12'd309,  12'd85,  
12'd224,  12'd227,  -12'd97,  12'd181,  12'd44,  12'd369,  -12'd168,  12'd376,  -12'd32,  12'd340,  12'd192,  12'd281,  12'd342,  12'd276,  -12'd65,  12'd50,  
-12'd130,  12'd207,  12'd265,  12'd158,  12'd42,  -12'd434,  12'd107,  12'd344,  12'd204,  -12'd294,  12'd293,  12'd230,  -12'd187,  -12'd84,  12'd187,  12'd415,  
12'd55,  12'd188,  -12'd0,  -12'd29,  -12'd144,  -12'd125,  12'd173,  -12'd47,  -12'd1,  -12'd62,  12'd70,  -12'd154,  -12'd82,  -12'd272,  12'd230,  -12'd86,  
-12'd215,  -12'd102,  12'd38,  -12'd234,  12'd181,  12'd8,  -12'd30,  12'd68,  12'd314,  12'd92,  12'd278,  12'd142,  -12'd317,  12'd37,  -12'd94,  12'd206,  
12'd5,  12'd431,  12'd123,  12'd150,  -12'd73,  -12'd32,  -12'd164,  12'd363,  12'd216,  -12'd149,  -12'd208,  -12'd170,  12'd186,  12'd457,  -12'd43,  -12'd142,  
12'd173,  -12'd258,  -12'd154,  12'd47,  12'd110,  -12'd44,  -12'd82,  12'd278,  
12'd189,  -12'd213,  -12'd89,  12'd22,  12'd133,  -12'd234,  -12'd200,  12'd209,  -12'd113,  12'd149,  -12'd509,  12'd114,  12'd49,  -12'd7,  12'd321,  -12'd371,  
12'd64,  -12'd53,  -12'd694,  -12'd107,  12'd280,  -12'd85,  -12'd154,  -12'd258,  -12'd283,  12'd121,  12'd33,  -12'd328,  -12'd114,  12'd403,  12'd157,  -12'd44,  
12'd233,  12'd356,  -12'd152,  12'd238,  12'd239,  12'd128,  -12'd263,  -12'd463,  12'd39,  12'd80,  12'd178,  -12'd701,  12'd366,  12'd27,  -12'd282,  -12'd288,  
-12'd276,  -12'd119,  12'd356,  -12'd469,  -12'd250,  12'd393,  -12'd104,  12'd165,  -12'd269,  -12'd16,  -12'd446,  12'd215,  -12'd194,  -12'd354,  12'd218,  12'd60,  
12'd38,  12'd138,  -12'd72,  -12'd229,  -12'd309,  12'd17,  12'd192,  -12'd198,  -12'd200,  12'd144,  12'd81,  12'd104,  12'd36,  12'd253,  12'd102,  12'd105,  
12'd133,  -12'd438,  -12'd243,  -12'd69,  12'd181,  12'd15,  12'd37,  12'd145,  -12'd496,  12'd100,  12'd120,  -12'd421,  -12'd24,  12'd333,  -12'd323,  12'd178,  
-12'd110,  12'd161,  -12'd72,  -12'd324,  12'd382,  -12'd44,  -12'd94,  12'd157,  -12'd48,  -12'd101,  -12'd252,  -12'd124,  -12'd215,  12'd5,  -12'd82,  12'd443,  
-12'd326,  12'd250,  12'd77,  12'd132,  -12'd250,  -12'd226,  12'd150,  -12'd50,  
12'd58,  -12'd204,  12'd261,  -12'd8,  12'd84,  12'd30,  12'd179,  -12'd57,  12'd106,  -12'd220,  12'd60,  12'd102,  -12'd361,  12'd55,  -12'd276,  -12'd269,  
12'd283,  12'd219,  12'd296,  12'd209,  -12'd196,  -12'd30,  12'd125,  -12'd41,  12'd316,  12'd141,  -12'd197,  -12'd125,  -12'd33,  12'd300,  -12'd313,  -12'd408,  
-12'd39,  12'd38,  12'd77,  12'd34,  -12'd236,  12'd281,  12'd34,  12'd349,  12'd133,  12'd75,  12'd230,  -12'd218,  -12'd207,  -12'd10,  12'd55,  12'd352,  
12'd4,  12'd161,  -12'd231,  12'd194,  -12'd502,  -12'd140,  12'd420,  -12'd266,  12'd118,  12'd206,  12'd12,  -12'd230,  12'd81,  -12'd280,  -12'd8,  -12'd177,  
-12'd133,  12'd149,  12'd31,  -12'd137,  12'd157,  12'd198,  12'd36,  12'd126,  -12'd73,  12'd18,  12'd2,  -12'd413,  12'd29,  12'd141,  -12'd32,  -12'd348,  
-12'd136,  -12'd267,  12'd314,  12'd442,  12'd292,  12'd191,  -12'd94,  -12'd293,  12'd301,  12'd313,  12'd238,  -12'd71,  -12'd381,  12'd453,  -12'd183,  12'd301,  
-12'd144,  -12'd111,  12'd268,  12'd249,  -12'd27,  12'd27,  12'd170,  12'd451,  -12'd116,  12'd19,  -12'd97,  12'd156,  12'd108,  -12'd420,  12'd433,  -12'd316,  
-12'd352,  -12'd256,  12'd51,  12'd69,  12'd183,  -12'd91,  -12'd74,  -12'd137,  
-12'd164,  12'd223,  -12'd477,  12'd276,  12'd110,  -12'd38,  -12'd31,  12'd40,  12'd57,  -12'd270,  -12'd433,  12'd241,  12'd446,  -12'd255,  -12'd173,  12'd1,  
-12'd44,  12'd16,  -12'd41,  -12'd21,  -12'd42,  12'd29,  12'd22,  -12'd55,  -12'd87,  -12'd415,  12'd207,  12'd57,  12'd59,  -12'd152,  12'd332,  -12'd377,  
-12'd106,  -12'd182,  -12'd94,  12'd165,  -12'd374,  12'd89,  12'd346,  -12'd73,  12'd210,  -12'd143,  -12'd329,  12'd74,  12'd119,  -12'd211,  12'd132,  12'd386,  
-12'd245,  -12'd573,  -12'd72,  -12'd166,  12'd257,  12'd272,  -12'd397,  -12'd45,  12'd286,  12'd115,  -12'd122,  -12'd389,  12'd505,  -12'd77,  12'd96,  -12'd84,  
12'd12,  12'd32,  -12'd192,  -12'd83,  12'd369,  -12'd116,  12'd123,  12'd389,  -12'd194,  12'd247,  -12'd76,  12'd389,  12'd195,  12'd361,  -12'd298,  -12'd91,  
12'd204,  12'd314,  -12'd384,  12'd182,  -12'd309,  12'd14,  12'd192,  12'd353,  12'd88,  12'd17,  12'd23,  12'd94,  -12'd92,  -12'd0,  -12'd180,  12'd416,  
-12'd86,  12'd36,  12'd233,  12'd331,  12'd43,  -12'd142,  12'd302,  12'd403,  -12'd157,  -12'd64,  12'd114,  12'd492,  12'd76,  -12'd17,  12'd221,  12'd141,  
-12'd38,  12'd440,  12'd257,  12'd52,  12'd384,  -12'd319,  12'd48,  -12'd74
};
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule


module bias_fc3_rom(
	input			clk,
	input							rstn,
	input	[`W_OUPTUT_BATCH:0]		aa,
	input							cena,
	output reg		[`WDP_BIAS*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	logic [0:`OUTPUT_BATCH_FC3-1][0:`OUTPUT_NUM_FC3-1][`WD_BIAS:0] weight	 = {
-24'd186531,  24'd166143,  -24'd211411,  -24'd80228,  -24'd155665,  24'd207658,  -24'd315652,  -24'd209780,  24'd326774,  24'd153726
	};

	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];	
endmodule




module wieght_fc3_rom(
	input			clk,
	input			rstn,
	input	[$clog2(`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3*`OUTPUT_BATCH_FC3)-1:0]	aa,
	input			cena,
	output reg		[`WDP*`OUTPUT_NUM_FC2*`OUTPUT_NUM_FC3 -1:0]	qa
	);
	
	
	//logic [0:`KERNEL_SIZE_CONV2*`KERNEL_SIZE_CONV2-1][0:`OUTPUT_NUM_CONV2-1][0:`OUTPUT_NUM_CONV1-1][31:0] weight	 = {
	logic [0:`OUTPUT_BATCH_FC3*`KERNEL_SIZEX_FC3*`KERNEL_SIZEY_FC3-1][0:`OUTPUT_NUM_FC3-1][0:`OUTPUT_NUM_FC2-1][`WD:0] weight	 = {
-12'd24,  12'd213,  -12'd32,  -12'd63,  12'd70,  12'd114,  12'd59,  -12'd54,  -12'd232,  -12'd180,  12'd510,  -12'd345,  -12'd113,  -12'd19,  -12'd256,  12'd204,  
12'd296,  12'd47,  -12'd48,  12'd521,  12'd648,  -12'd489,  -12'd343,  -12'd44,  -12'd403,  12'd327,  12'd125,  -12'd38,  -12'd186,  12'd249,  12'd85,  12'd308,  
-12'd293,  -12'd494,  -12'd171,  -12'd471,  -12'd131,  12'd175,  12'd126,  -12'd129,  12'd193,  -12'd35,  12'd365,  -12'd170,  -12'd438,  12'd88,  -12'd91,  12'd82,  
-12'd511,  -12'd66,  12'd298,  12'd80,  12'd511,  -12'd181,  -12'd315,  12'd289,  -12'd188,  12'd517,  12'd1,  -12'd65,  -12'd117,  -12'd120,  12'd91,  -12'd289,  
12'd428,  -12'd457,  -12'd121,  -12'd87,  -12'd232,  -12'd255,  -12'd19,  -12'd610,  -12'd28,  -12'd136,  -12'd232,  12'd75,  12'd48,  -12'd178,  12'd300,  -12'd98,  
-12'd118,  -12'd292,  12'd388,  -12'd261,  
12'd285,  -12'd427,  12'd83,  -12'd198,  -12'd28,  12'd105,  12'd214,  -12'd162,  -12'd36,  -12'd261,  -12'd480,  12'd239,  12'd29,  12'd344,  12'd126,  12'd124,  
-12'd289,  12'd262,  -12'd258,  -12'd198,  12'd445,  -12'd137,  -12'd13,  12'd35,  -12'd437,  -12'd50,  -12'd84,  12'd329,  12'd248,  -12'd51,  12'd337,  -12'd113,  
12'd4,  -12'd268,  -12'd2,  12'd402,  -12'd225,  -12'd246,  -12'd127,  -12'd394,  12'd304,  -12'd193,  -12'd574,  -12'd434,  12'd280,  12'd196,  -12'd1,  12'd196,  
-12'd213,  12'd346,  -12'd489,  -12'd216,  -12'd68,  12'd200,  12'd522,  -12'd247,  -12'd130,  -12'd158,  -12'd578,  12'd503,  -12'd255,  12'd60,  -12'd356,  -12'd113,  
12'd393,  -12'd236,  12'd128,  12'd559,  12'd184,  -12'd366,  -12'd250,  12'd311,  12'd232,  12'd65,  -12'd401,  -12'd225,  -12'd23,  -12'd422,  -12'd351,  12'd128,  
12'd212,  -12'd503,  12'd502,  -12'd78,  
-12'd353,  -12'd359,  12'd229,  -12'd48,  12'd483,  12'd197,  -12'd198,  12'd47,  12'd135,  -12'd192,  12'd233,  12'd424,  12'd78,  -12'd333,  -12'd122,  -12'd159,  
-12'd69,  -12'd630,  -12'd329,  12'd209,  12'd399,  12'd54,  -12'd162,  -12'd338,  12'd26,  -12'd107,  -12'd43,  -12'd123,  -12'd193,  12'd373,  -12'd663,  -12'd27,  
-12'd617,  -12'd121,  12'd26,  -12'd329,  12'd85,  12'd288,  12'd98,  12'd452,  -12'd27,  -12'd94,  12'd94,  -12'd204,  12'd28,  -12'd50,  12'd231,  12'd205,  
12'd262,  12'd299,  -12'd561,  -12'd434,  -12'd128,  -12'd148,  -12'd212,  -12'd171,  12'd83,  12'd301,  12'd7,  12'd106,  -12'd35,  -12'd421,  -12'd31,  12'd320,  
12'd146,  -12'd326,  12'd104,  -12'd242,  -12'd140,  12'd158,  12'd149,  12'd88,  -12'd286,  12'd176,  -12'd235,  12'd41,  -12'd94,  12'd425,  12'd108,  -12'd322,  
12'd473,  -12'd101,  -12'd26,  -12'd243,  
-12'd2,  -12'd223,  12'd33,  -12'd479,  12'd276,  12'd42,  -12'd246,  -12'd211,  12'd86,  -12'd150,  -12'd321,  -12'd250,  12'd475,  -12'd286,  -12'd283,  12'd89,  
-12'd279,  12'd141,  -12'd191,  12'd378,  -12'd631,  -12'd253,  -12'd278,  -12'd375,  -12'd29,  12'd102,  -12'd301,  12'd94,  -12'd330,  12'd240,  -12'd65,  -12'd94,  
12'd34,  12'd127,  -12'd272,  12'd252,  12'd145,  -12'd224,  -12'd87,  12'd248,  -12'd215,  -12'd110,  12'd333,  12'd161,  12'd282,  -12'd394,  -12'd148,  -12'd242,  
12'd302,  -12'd472,  12'd50,  12'd348,  -12'd330,  -12'd9,  -12'd117,  -12'd191,  -12'd202,  -12'd174,  12'd229,  12'd16,  12'd44,  12'd71,  -12'd38,  12'd114,  
-12'd383,  12'd648,  -12'd65,  12'd171,  12'd11,  12'd10,  -12'd396,  12'd307,  -12'd465,  12'd205,  -12'd142,  12'd4,  12'd288,  12'd31,  12'd2,  -12'd119,  
-12'd443,  -12'd116,  12'd70,  12'd511,  
-12'd296,  12'd328,  12'd15,  12'd113,  -12'd322,  12'd193,  12'd519,  12'd277,  -12'd406,  -12'd4,  -12'd145,  -12'd246,  -12'd165,  12'd367,  12'd208,  -12'd373,  
12'd358,  -12'd206,  -12'd488,  -12'd74,  -12'd331,  12'd174,  -12'd50,  -12'd508,  12'd211,  -12'd103,  -12'd759,  -12'd118,  12'd422,  12'd156,  -12'd394,  -12'd316,  
12'd7,  -12'd418,  -12'd100,  12'd36,  -12'd335,  12'd221,  12'd267,  -12'd443,  12'd2,  -12'd128,  12'd26,  12'd427,  12'd104,  12'd255,  -12'd74,  12'd93,  
12'd199,  -12'd133,  12'd221,  -12'd210,  12'd245,  12'd2,  -12'd176,  -12'd86,  -12'd60,  12'd95,  -12'd177,  12'd401,  -12'd19,  -12'd72,  -12'd311,  12'd294,  
12'd104,  -12'd401,  12'd39,  12'd397,  -12'd490,  -12'd241,  12'd339,  -12'd226,  -12'd445,  -12'd356,  12'd240,  12'd350,  -12'd410,  12'd231,  -12'd423,  12'd321,  
-12'd320,  12'd232,  -12'd269,  -12'd317,  
12'd556,  12'd279,  -12'd369,  -12'd369,  12'd506,  -12'd313,  -12'd384,  12'd126,  12'd294,  12'd301,  12'd115,  12'd511,  -12'd347,  -12'd296,  12'd44,  -12'd180,  
12'd147,  12'd376,  12'd213,  12'd206,  -12'd307,  12'd160,  -12'd231,  12'd336,  12'd313,  12'd174,  12'd225,  12'd50,  -12'd171,  12'd14,  12'd112,  -12'd160,  
-12'd6,  -12'd59,  12'd142,  12'd537,  -12'd305,  -12'd564,  -12'd455,  12'd129,  12'd204,  12'd16,  -12'd338,  -12'd280,  -12'd332,  -12'd223,  -12'd158,  12'd0,  
12'd309,  12'd338,  12'd43,  12'd308,  12'd119,  -12'd452,  -12'd514,  12'd128,  -12'd172,  -12'd108,  12'd136,  -12'd349,  12'd1,  12'd13,  12'd23,  -12'd383,  
-12'd22,  -12'd90,  12'd341,  12'd89,  -12'd43,  -12'd225,  -12'd166,  -12'd35,  12'd509,  -12'd42,  12'd284,  12'd129,  12'd127,  -12'd96,  12'd12,  12'd271,  
-12'd375,  12'd168,  -12'd359,  12'd81,  
12'd463,  -12'd252,  -12'd56,  -12'd14,  -12'd23,  -12'd326,  -12'd57,  12'd274,  12'd103,  12'd278,  -12'd196,  -12'd281,  -12'd757,  -12'd43,  -12'd305,  -12'd293,  
12'd285,  -12'd109,  -12'd380,  -12'd260,  12'd83,  12'd88,  -12'd362,  -12'd178,  12'd188,  -12'd153,  -12'd14,  12'd10,  -12'd424,  12'd49,  12'd277,  12'd177,  
-12'd173,  12'd435,  -12'd31,  -12'd130,  -12'd371,  -12'd320,  12'd201,  -12'd204,  -12'd159,  -12'd367,  12'd542,  -12'd452,  12'd37,  -12'd139,  12'd196,  -12'd30,  
-12'd129,  -12'd391,  12'd266,  -12'd239,  12'd24,  12'd226,  12'd67,  12'd192,  -12'd0,  12'd100,  12'd156,  -12'd6,  12'd161,  -12'd358,  12'd164,  -12'd466,  
12'd139,  12'd231,  -12'd64,  12'd25,  -12'd26,  12'd103,  12'd159,  -12'd258,  12'd244,  -12'd176,  12'd111,  -12'd355,  -12'd270,  12'd162,  -12'd250,  12'd62,  
12'd132,  12'd201,  -12'd203,  -12'd612,  
-12'd353,  -12'd81,  12'd172,  -12'd674,  -12'd275,  12'd175,  -12'd565,  -12'd172,  -12'd219,  -12'd189,  -12'd564,  12'd112,  12'd84,  12'd157,  -12'd239,  12'd33,  
12'd225,  -12'd22,  -12'd232,  -12'd151,  -12'd133,  -12'd170,  -12'd213,  -12'd199,  -12'd107,  -12'd44,  -12'd53,  -12'd189,  12'd453,  -12'd98,  12'd151,  -12'd22,  
12'd10,  -12'd88,  12'd558,  -12'd178,  12'd64,  12'd419,  -12'd338,  -12'd125,  -12'd139,  12'd82,  -12'd565,  -12'd15,  12'd407,  12'd415,  -12'd169,  -12'd78,  
12'd61,  12'd110,  12'd166,  -12'd385,  12'd190,  12'd66,  12'd37,  -12'd282,  12'd156,  -12'd656,  -12'd382,  12'd240,  -12'd49,  12'd336,  -12'd252,  -12'd245,  
-12'd58,  12'd522,  12'd15,  -12'd593,  12'd366,  -12'd162,  12'd46,  12'd18,  12'd58,  -12'd58,  12'd162,  12'd68,  12'd258,  12'd206,  12'd267,  -12'd20,  
12'd174,  -12'd381,  12'd87,  12'd2,  
12'd25,  12'd262,  12'd193,  -12'd55,  -12'd9,  -12'd14,  12'd3,  -12'd208,  -12'd68,  12'd522,  -12'd423,  -12'd502,  12'd60,  -12'd393,  -12'd20,  12'd67,  
12'd117,  12'd154,  12'd244,  12'd64,  12'd34,  12'd295,  -12'd49,  -12'd190,  12'd30,  -12'd232,  -12'd375,  12'd42,  -12'd284,  -12'd200,  -12'd555,  -12'd240,  
-12'd367,  12'd231,  -12'd202,  12'd223,  12'd64,  12'd37,  -12'd61,  12'd143,  -12'd38,  12'd61,  -12'd254,  12'd470,  -12'd352,  12'd325,  12'd62,  12'd71,  
-12'd336,  -12'd473,  -12'd319,  12'd290,  12'd264,  12'd260,  12'd161,  12'd130,  -12'd72,  -12'd303,  12'd84,  -12'd317,  12'd347,  -12'd314,  12'd284,  -12'd0,  
12'd238,  12'd302,  -12'd310,  -12'd192,  12'd13,  -12'd442,  -12'd390,  12'd4,  12'd210,  12'd23,  12'd135,  -12'd463,  -12'd313,  12'd39,  12'd84,  -12'd479,  
12'd316,  12'd449,  -12'd14,  -12'd87,  
12'd98,  12'd126,  12'd186,  12'd100,  12'd177,  -12'd216,  12'd168,  12'd147,  -12'd196,  -12'd275,  12'd162,  12'd207,  12'd311,  12'd347,  12'd202,  12'd106,  
-12'd401,  -12'd33,  -12'd112,  -12'd177,  -12'd5,  -12'd189,  12'd269,  12'd66,  12'd295,  -12'd101,  12'd109,  -12'd146,  12'd147,  -12'd572,  -12'd280,  -12'd120,  
12'd51,  -12'd364,  12'd101,  -12'd44,  -12'd205,  12'd408,  12'd151,  12'd316,  12'd353,  12'd319,  -12'd143,  12'd67,  12'd184,  -12'd62,  12'd74,  -12'd34,  
-12'd572,  -12'd183,  -12'd48,  12'd204,  12'd221,  -12'd41,  -12'd660,  -12'd33,  -12'd66,  12'd277,  12'd170,  -12'd485,  12'd47,  12'd236,  12'd574,  12'd285,  
-12'd120,  -12'd738,  12'd135,  12'd61,  -12'd6,  12'd387,  12'd329,  12'd255,  -12'd142,  -12'd659,  12'd325,  -12'd419,  -12'd60,  -12'd462,  -12'd332,  12'd110,  
-12'd407,  -12'd332,  -12'd142,  -12'd11
	};
	
	always @(`CLK_RST_EDGE)
		if (`RST)			qa <= 0;
		else if (!cena)		qa <= weight[aa];
endmodule

